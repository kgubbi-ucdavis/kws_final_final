VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CNN_Accelerator_Top
  CLASS BLOCK ;
  FOREIGN CNN_Accelerator_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 820.000 BY 800.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END done
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END reset
  PIN serial_line_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 796.000 341.690 800.000 ;
    END
  END serial_line_data[0]
  PIN serial_line_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 204.790 796.000 205.070 800.000 ;
    END
  END serial_line_data[1]
  PIN serial_line_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 68.170 796.000 68.450 800.000 ;
    END
  END serial_line_data[2]
  PIN serial_line_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 816.000 731.720 820.000 732.320 ;
    END
  END serial_line_data[3]
  PIN serial_line_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 816.000 598.440 820.000 599.040 ;
    END
  END serial_line_data[4]
  PIN serial_line_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 816.000 465.160 820.000 465.760 ;
    END
  END serial_line_data[5]
  PIN serial_line_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 816.000 331.880 820.000 332.480 ;
    END
  END serial_line_data[6]
  PIN serial_line_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 816.000 198.600 820.000 199.200 ;
    END
  END serial_line_data[7]
  PIN serial_line_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 478.030 796.000 478.310 800.000 ;
    END
  END serial_line_valid
  PIN serial_result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END serial_result[0]
  PIN serial_result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END serial_result[1]
  PIN serial_result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END serial_result[2]
  PIN serial_result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END serial_result[3]
  PIN serial_result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END serial_result[4]
  PIN serial_result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END serial_result[5]
  PIN serial_result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 751.270 796.000 751.550 800.000 ;
    END
  END serial_result[6]
  PIN serial_result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 614.650 796.000 614.930 800.000 ;
    END
  END serial_result[7]
  PIN serial_result_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END serial_result_valid
  PIN serial_weight_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END serial_weight_data[0]
  PIN serial_weight_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END serial_weight_data[1]
  PIN serial_weight_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END serial_weight_data[2]
  PIN serial_weight_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END serial_weight_data[3]
  PIN serial_weight_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END serial_weight_data[4]
  PIN serial_weight_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END serial_weight_data[5]
  PIN serial_weight_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END serial_weight_data[6]
  PIN serial_weight_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END serial_weight_data[7]
  PIN serial_weight_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 816.000 65.320 820.000 65.920 ;
    END
  END serial_weight_valid
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 814.200 788.885 ;
      LAYER met1 ;
        RECT 5.520 10.640 814.200 789.040 ;
      LAYER met2 ;
        RECT 6.530 795.720 67.890 796.000 ;
        RECT 68.730 795.720 204.510 796.000 ;
        RECT 205.350 795.720 341.130 796.000 ;
        RECT 341.970 795.720 477.750 796.000 ;
        RECT 478.590 795.720 614.370 796.000 ;
        RECT 615.210 795.720 750.990 796.000 ;
        RECT 751.830 795.720 814.110 796.000 ;
        RECT 6.530 4.280 814.110 795.720 ;
        RECT 6.530 3.670 36.610 4.280 ;
        RECT 37.450 3.670 111.130 4.280 ;
        RECT 111.970 3.670 185.650 4.280 ;
        RECT 186.490 3.670 260.170 4.280 ;
        RECT 261.010 3.670 334.690 4.280 ;
        RECT 335.530 3.670 409.210 4.280 ;
        RECT 410.050 3.670 483.730 4.280 ;
        RECT 484.570 3.670 558.250 4.280 ;
        RECT 559.090 3.670 632.770 4.280 ;
        RECT 633.610 3.670 707.290 4.280 ;
        RECT 708.130 3.670 781.810 4.280 ;
        RECT 782.650 3.670 814.110 4.280 ;
      LAYER met3 ;
        RECT 4.000 747.680 816.000 788.965 ;
        RECT 4.400 746.280 816.000 747.680 ;
        RECT 4.000 732.720 816.000 746.280 ;
        RECT 4.000 731.320 815.600 732.720 ;
        RECT 4.000 648.400 816.000 731.320 ;
        RECT 4.400 647.000 816.000 648.400 ;
        RECT 4.000 599.440 816.000 647.000 ;
        RECT 4.000 598.040 815.600 599.440 ;
        RECT 4.000 549.120 816.000 598.040 ;
        RECT 4.400 547.720 816.000 549.120 ;
        RECT 4.000 466.160 816.000 547.720 ;
        RECT 4.000 464.760 815.600 466.160 ;
        RECT 4.000 449.840 816.000 464.760 ;
        RECT 4.400 448.440 816.000 449.840 ;
        RECT 4.000 350.560 816.000 448.440 ;
        RECT 4.400 349.160 816.000 350.560 ;
        RECT 4.000 332.880 816.000 349.160 ;
        RECT 4.000 331.480 815.600 332.880 ;
        RECT 4.000 251.280 816.000 331.480 ;
        RECT 4.400 249.880 816.000 251.280 ;
        RECT 4.000 199.600 816.000 249.880 ;
        RECT 4.000 198.200 815.600 199.600 ;
        RECT 4.000 152.000 816.000 198.200 ;
        RECT 4.400 150.600 816.000 152.000 ;
        RECT 4.000 66.320 816.000 150.600 ;
        RECT 4.000 64.920 815.600 66.320 ;
        RECT 4.000 52.720 816.000 64.920 ;
        RECT 4.400 51.320 816.000 52.720 ;
        RECT 4.000 10.715 816.000 51.320 ;
      LAYER met4 ;
        RECT 230.295 11.735 251.040 713.825 ;
        RECT 253.440 11.735 327.840 713.825 ;
        RECT 330.240 11.735 404.640 713.825 ;
        RECT 407.040 11.735 481.440 713.825 ;
        RECT 483.840 11.735 558.240 713.825 ;
        RECT 560.640 11.735 563.665 713.825 ;
  END
END CNN_Accelerator_Top
END LIBRARY


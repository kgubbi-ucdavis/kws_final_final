VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CNN_Accelerator_Top
  CLASS BLOCK ;
  FOREIGN CNN_Accelerator_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 820.000 BY 800.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END done
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END reset
  PIN serial_line_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END serial_line_data[0]
  PIN serial_line_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END serial_line_data[1]
  PIN serial_line_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END serial_line_data[2]
  PIN serial_line_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END serial_line_data[3]
  PIN serial_line_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END serial_line_data[4]
  PIN serial_line_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END serial_line_data[5]
  PIN serial_line_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END serial_line_data[6]
  PIN serial_line_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END serial_line_data[7]
  PIN serial_line_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END serial_line_valid
  PIN serial_result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END serial_result[0]
  PIN serial_result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END serial_result[1]
  PIN serial_result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END serial_result[2]
  PIN serial_result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END serial_result[3]
  PIN serial_result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END serial_result[4]
  PIN serial_result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END serial_result[5]
  PIN serial_result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 4.000 ;
    END
  END serial_result[6]
  PIN serial_result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END serial_result[7]
  PIN serial_result_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 776.570 0.000 776.850 4.000 ;
    END
  END serial_result_valid
  PIN serial_weight_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END serial_weight_data[0]
  PIN serial_weight_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END serial_weight_data[1]
  PIN serial_weight_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END serial_weight_data[2]
  PIN serial_weight_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END serial_weight_data[3]
  PIN serial_weight_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END serial_weight_data[4]
  PIN serial_weight_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END serial_weight_data[5]
  PIN serial_weight_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END serial_weight_data[6]
  PIN serial_weight_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END serial_weight_data[7]
  PIN serial_weight_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END serial_weight_valid
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 784.665 814.390 787.495 ;
        RECT 5.330 779.225 814.390 782.055 ;
        RECT 5.330 773.785 814.390 776.615 ;
        RECT 5.330 768.345 814.390 771.175 ;
        RECT 5.330 762.905 814.390 765.735 ;
        RECT 5.330 757.465 814.390 760.295 ;
        RECT 5.330 752.025 814.390 754.855 ;
        RECT 5.330 746.585 814.390 749.415 ;
        RECT 5.330 741.145 814.390 743.975 ;
        RECT 5.330 735.705 814.390 738.535 ;
        RECT 5.330 730.265 814.390 733.095 ;
        RECT 5.330 724.825 814.390 727.655 ;
        RECT 5.330 719.385 814.390 722.215 ;
        RECT 5.330 713.945 814.390 716.775 ;
        RECT 5.330 708.505 814.390 711.335 ;
        RECT 5.330 703.065 814.390 705.895 ;
        RECT 5.330 697.625 814.390 700.455 ;
        RECT 5.330 692.185 814.390 695.015 ;
        RECT 5.330 686.745 814.390 689.575 ;
        RECT 5.330 681.305 814.390 684.135 ;
        RECT 5.330 675.865 814.390 678.695 ;
        RECT 5.330 670.425 814.390 673.255 ;
        RECT 5.330 664.985 814.390 667.815 ;
        RECT 5.330 659.545 814.390 662.375 ;
        RECT 5.330 654.105 814.390 656.935 ;
        RECT 5.330 648.665 814.390 651.495 ;
        RECT 5.330 643.225 814.390 646.055 ;
        RECT 5.330 637.785 814.390 640.615 ;
        RECT 5.330 632.345 814.390 635.175 ;
        RECT 5.330 626.905 814.390 629.735 ;
        RECT 5.330 621.465 814.390 624.295 ;
        RECT 5.330 616.025 814.390 618.855 ;
        RECT 5.330 610.585 814.390 613.415 ;
        RECT 5.330 605.145 814.390 607.975 ;
        RECT 5.330 599.705 814.390 602.535 ;
        RECT 5.330 594.265 814.390 597.095 ;
        RECT 5.330 588.825 814.390 591.655 ;
        RECT 5.330 583.385 814.390 586.215 ;
        RECT 5.330 577.945 814.390 580.775 ;
        RECT 5.330 572.505 814.390 575.335 ;
        RECT 5.330 567.065 814.390 569.895 ;
        RECT 5.330 561.625 814.390 564.455 ;
        RECT 5.330 556.185 814.390 559.015 ;
        RECT 5.330 550.745 814.390 553.575 ;
        RECT 5.330 545.305 814.390 548.135 ;
        RECT 5.330 539.865 814.390 542.695 ;
        RECT 5.330 534.425 814.390 537.255 ;
        RECT 5.330 528.985 814.390 531.815 ;
        RECT 5.330 523.545 814.390 526.375 ;
        RECT 5.330 518.105 814.390 520.935 ;
        RECT 5.330 512.665 814.390 515.495 ;
        RECT 5.330 507.225 814.390 510.055 ;
        RECT 5.330 501.785 814.390 504.615 ;
        RECT 5.330 496.345 814.390 499.175 ;
        RECT 5.330 490.905 814.390 493.735 ;
        RECT 5.330 485.465 814.390 488.295 ;
        RECT 5.330 480.025 814.390 482.855 ;
        RECT 5.330 474.585 814.390 477.415 ;
        RECT 5.330 469.145 814.390 471.975 ;
        RECT 5.330 463.705 814.390 466.535 ;
        RECT 5.330 458.265 814.390 461.095 ;
        RECT 5.330 452.825 814.390 455.655 ;
        RECT 5.330 447.385 814.390 450.215 ;
        RECT 5.330 441.945 814.390 444.775 ;
        RECT 5.330 436.505 814.390 439.335 ;
        RECT 5.330 431.065 814.390 433.895 ;
        RECT 5.330 425.625 814.390 428.455 ;
        RECT 5.330 420.185 814.390 423.015 ;
        RECT 5.330 414.745 814.390 417.575 ;
        RECT 5.330 409.305 814.390 412.135 ;
        RECT 5.330 403.865 814.390 406.695 ;
        RECT 5.330 398.425 814.390 401.255 ;
        RECT 5.330 392.985 814.390 395.815 ;
        RECT 5.330 387.545 814.390 390.375 ;
        RECT 5.330 382.105 814.390 384.935 ;
        RECT 5.330 376.665 814.390 379.495 ;
        RECT 5.330 371.225 814.390 374.055 ;
        RECT 5.330 365.785 814.390 368.615 ;
        RECT 5.330 360.345 814.390 363.175 ;
        RECT 5.330 354.905 814.390 357.735 ;
        RECT 5.330 349.465 814.390 352.295 ;
        RECT 5.330 344.025 814.390 346.855 ;
        RECT 5.330 338.585 814.390 341.415 ;
        RECT 5.330 333.145 814.390 335.975 ;
        RECT 5.330 327.705 814.390 330.535 ;
        RECT 5.330 322.265 814.390 325.095 ;
        RECT 5.330 316.825 814.390 319.655 ;
        RECT 5.330 311.385 814.390 314.215 ;
        RECT 5.330 305.945 814.390 308.775 ;
        RECT 5.330 300.505 814.390 303.335 ;
        RECT 5.330 295.065 814.390 297.895 ;
        RECT 5.330 289.625 814.390 292.455 ;
        RECT 5.330 284.185 814.390 287.015 ;
        RECT 5.330 278.745 814.390 281.575 ;
        RECT 5.330 273.305 814.390 276.135 ;
        RECT 5.330 267.865 814.390 270.695 ;
        RECT 5.330 262.425 814.390 265.255 ;
        RECT 5.330 256.985 814.390 259.815 ;
        RECT 5.330 251.545 814.390 254.375 ;
        RECT 5.330 246.105 814.390 248.935 ;
        RECT 5.330 240.665 814.390 243.495 ;
        RECT 5.330 235.225 814.390 238.055 ;
        RECT 5.330 229.785 814.390 232.615 ;
        RECT 5.330 224.345 814.390 227.175 ;
        RECT 5.330 218.905 814.390 221.735 ;
        RECT 5.330 213.465 814.390 216.295 ;
        RECT 5.330 208.025 814.390 210.855 ;
        RECT 5.330 202.585 814.390 205.415 ;
        RECT 5.330 197.145 814.390 199.975 ;
        RECT 5.330 191.705 814.390 194.535 ;
        RECT 5.330 186.265 814.390 189.095 ;
        RECT 5.330 180.825 814.390 183.655 ;
        RECT 5.330 175.385 814.390 178.215 ;
        RECT 5.330 169.945 814.390 172.775 ;
        RECT 5.330 164.505 814.390 167.335 ;
        RECT 5.330 159.065 814.390 161.895 ;
        RECT 5.330 153.625 814.390 156.455 ;
        RECT 5.330 148.185 814.390 151.015 ;
        RECT 5.330 142.745 814.390 145.575 ;
        RECT 5.330 137.305 814.390 140.135 ;
        RECT 5.330 131.865 814.390 134.695 ;
        RECT 5.330 126.425 814.390 129.255 ;
        RECT 5.330 120.985 814.390 123.815 ;
        RECT 5.330 115.545 814.390 118.375 ;
        RECT 5.330 110.105 814.390 112.935 ;
        RECT 5.330 104.665 814.390 107.495 ;
        RECT 5.330 99.225 814.390 102.055 ;
        RECT 5.330 93.785 814.390 96.615 ;
        RECT 5.330 88.345 814.390 91.175 ;
        RECT 5.330 82.905 814.390 85.735 ;
        RECT 5.330 77.465 814.390 80.295 ;
        RECT 5.330 72.025 814.390 74.855 ;
        RECT 5.330 66.585 814.390 69.415 ;
        RECT 5.330 61.145 814.390 63.975 ;
        RECT 5.330 55.705 814.390 58.535 ;
        RECT 5.330 50.265 814.390 53.095 ;
        RECT 5.330 44.825 814.390 47.655 ;
        RECT 5.330 39.385 814.390 42.215 ;
        RECT 5.330 33.945 814.390 36.775 ;
        RECT 5.330 28.505 814.390 31.335 ;
        RECT 5.330 23.065 814.390 25.895 ;
        RECT 5.330 17.625 814.390 20.455 ;
        RECT 5.330 12.185 814.390 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 814.200 788.885 ;
      LAYER met1 ;
        RECT 5.520 8.880 814.200 789.040 ;
      LAYER met2 ;
        RECT 16.200 4.280 805.360 788.985 ;
        RECT 16.750 3.670 42.130 4.280 ;
        RECT 42.970 3.670 68.350 4.280 ;
        RECT 69.190 3.670 94.570 4.280 ;
        RECT 95.410 3.670 120.790 4.280 ;
        RECT 121.630 3.670 147.010 4.280 ;
        RECT 147.850 3.670 173.230 4.280 ;
        RECT 174.070 3.670 199.450 4.280 ;
        RECT 200.290 3.670 225.670 4.280 ;
        RECT 226.510 3.670 251.890 4.280 ;
        RECT 252.730 3.670 278.110 4.280 ;
        RECT 278.950 3.670 304.330 4.280 ;
        RECT 305.170 3.670 330.550 4.280 ;
        RECT 331.390 3.670 356.770 4.280 ;
        RECT 357.610 3.670 382.990 4.280 ;
        RECT 383.830 3.670 409.210 4.280 ;
        RECT 410.050 3.670 435.430 4.280 ;
        RECT 436.270 3.670 461.650 4.280 ;
        RECT 462.490 3.670 487.870 4.280 ;
        RECT 488.710 3.670 514.090 4.280 ;
        RECT 514.930 3.670 540.310 4.280 ;
        RECT 541.150 3.670 566.530 4.280 ;
        RECT 567.370 3.670 592.750 4.280 ;
        RECT 593.590 3.670 618.970 4.280 ;
        RECT 619.810 3.670 645.190 4.280 ;
        RECT 646.030 3.670 671.410 4.280 ;
        RECT 672.250 3.670 697.630 4.280 ;
        RECT 698.470 3.670 723.850 4.280 ;
        RECT 724.690 3.670 750.070 4.280 ;
        RECT 750.910 3.670 776.290 4.280 ;
        RECT 777.130 3.670 802.510 4.280 ;
        RECT 803.350 3.670 805.360 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 790.630 788.965 ;
      LAYER met4 ;
        RECT 229.375 17.175 251.040 409.185 ;
        RECT 253.440 17.175 327.840 409.185 ;
        RECT 330.240 17.175 404.640 409.185 ;
        RECT 407.040 17.175 481.440 409.185 ;
        RECT 483.840 17.175 558.240 409.185 ;
        RECT 560.640 17.175 569.185 409.185 ;
  END
END CNN_Accelerator_Top
END LIBRARY


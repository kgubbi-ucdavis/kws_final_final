magic
tech sky130A
magscale 1 2
timestamp 1717390112
<< nwell >>
rect 1066 156933 162878 157499
rect 1066 155845 162878 156411
rect 1066 154757 162878 155323
rect 1066 153669 162878 154235
rect 1066 152581 162878 153147
rect 1066 151493 162878 152059
rect 1066 150405 162878 150971
rect 1066 149317 162878 149883
rect 1066 148229 162878 148795
rect 1066 147141 162878 147707
rect 1066 146053 162878 146619
rect 1066 144965 162878 145531
rect 1066 143877 162878 144443
rect 1066 142789 162878 143355
rect 1066 141701 162878 142267
rect 1066 140613 162878 141179
rect 1066 139525 162878 140091
rect 1066 138437 162878 139003
rect 1066 137349 162878 137915
rect 1066 136261 162878 136827
rect 1066 135173 162878 135739
rect 1066 134085 162878 134651
rect 1066 132997 162878 133563
rect 1066 131909 162878 132475
rect 1066 130821 162878 131387
rect 1066 129733 162878 130299
rect 1066 128645 162878 129211
rect 1066 127557 162878 128123
rect 1066 126469 162878 127035
rect 1066 125381 162878 125947
rect 1066 124293 162878 124859
rect 1066 123205 162878 123771
rect 1066 122117 162878 122683
rect 1066 121029 162878 121595
rect 1066 119941 162878 120507
rect 1066 118853 162878 119419
rect 1066 117765 162878 118331
rect 1066 116677 162878 117243
rect 1066 115589 162878 116155
rect 1066 114501 162878 115067
rect 1066 113413 162878 113979
rect 1066 112325 162878 112891
rect 1066 111237 162878 111803
rect 1066 110149 162878 110715
rect 1066 109061 162878 109627
rect 1066 107973 162878 108539
rect 1066 106885 162878 107451
rect 1066 105797 162878 106363
rect 1066 104709 162878 105275
rect 1066 103621 162878 104187
rect 1066 102533 162878 103099
rect 1066 101445 162878 102011
rect 1066 100357 162878 100923
rect 1066 99269 162878 99835
rect 1066 98181 162878 98747
rect 1066 97093 162878 97659
rect 1066 96005 162878 96571
rect 1066 94917 162878 95483
rect 1066 93829 162878 94395
rect 1066 92741 162878 93307
rect 1066 91653 162878 92219
rect 1066 90565 162878 91131
rect 1066 89477 162878 90043
rect 1066 88389 162878 88955
rect 1066 87301 162878 87867
rect 1066 86213 162878 86779
rect 1066 85125 162878 85691
rect 1066 84037 162878 84603
rect 1066 82949 162878 83515
rect 1066 81861 162878 82427
rect 1066 80773 162878 81339
rect 1066 79685 162878 80251
rect 1066 78597 162878 79163
rect 1066 77509 162878 78075
rect 1066 76421 162878 76987
rect 1066 75333 162878 75899
rect 1066 74245 162878 74811
rect 1066 73157 162878 73723
rect 1066 72069 162878 72635
rect 1066 70981 162878 71547
rect 1066 69893 162878 70459
rect 1066 68805 162878 69371
rect 1066 67717 162878 68283
rect 1066 66629 162878 67195
rect 1066 65541 162878 66107
rect 1066 64453 162878 65019
rect 1066 63365 162878 63931
rect 1066 62277 162878 62843
rect 1066 61189 162878 61755
rect 1066 60101 162878 60667
rect 1066 59013 162878 59579
rect 1066 57925 162878 58491
rect 1066 56837 162878 57403
rect 1066 55749 162878 56315
rect 1066 54661 162878 55227
rect 1066 53573 162878 54139
rect 1066 52485 162878 53051
rect 1066 51397 162878 51963
rect 1066 50309 162878 50875
rect 1066 49221 162878 49787
rect 1066 48133 162878 48699
rect 1066 47045 162878 47611
rect 1066 45957 162878 46523
rect 1066 44869 162878 45435
rect 1066 43781 162878 44347
rect 1066 42693 162878 43259
rect 1066 41605 162878 42171
rect 1066 40517 162878 41083
rect 1066 39429 162878 39995
rect 1066 38341 162878 38907
rect 1066 37253 162878 37819
rect 1066 36165 162878 36731
rect 1066 35077 162878 35643
rect 1066 33989 162878 34555
rect 1066 32901 162878 33467
rect 1066 31813 162878 32379
rect 1066 30725 162878 31291
rect 1066 29637 162878 30203
rect 1066 28549 162878 29115
rect 1066 27461 162878 28027
rect 1066 26373 162878 26939
rect 1066 25285 162878 25851
rect 1066 24197 162878 24763
rect 1066 23109 162878 23675
rect 1066 22021 162878 22587
rect 1066 20933 162878 21499
rect 1066 19845 162878 20411
rect 1066 18757 162878 19323
rect 1066 17669 162878 18235
rect 1066 16581 162878 17147
rect 1066 15493 162878 16059
rect 1066 14405 162878 14971
rect 1066 13317 162878 13883
rect 1066 12229 162878 12795
rect 1066 11141 162878 11707
rect 1066 10053 162878 10619
rect 1066 8965 162878 9531
rect 1066 7877 162878 8443
rect 1066 6789 162878 7355
rect 1066 5701 162878 6267
rect 1066 4613 162878 5179
rect 1066 3525 162878 4091
rect 1066 2437 162878 3003
<< obsli1 >>
rect 1104 2159 162840 157777
<< obsm1 >>
rect 1104 1776 162840 157808
<< metal2 >>
rect 3238 0 3294 800
rect 8482 0 8538 800
rect 13726 0 13782 800
rect 18970 0 19026 800
rect 24214 0 24270 800
rect 29458 0 29514 800
rect 34702 0 34758 800
rect 39946 0 40002 800
rect 45190 0 45246 800
rect 50434 0 50490 800
rect 55678 0 55734 800
rect 60922 0 60978 800
rect 66166 0 66222 800
rect 71410 0 71466 800
rect 76654 0 76710 800
rect 81898 0 81954 800
rect 87142 0 87198 800
rect 92386 0 92442 800
rect 97630 0 97686 800
rect 102874 0 102930 800
rect 108118 0 108174 800
rect 113362 0 113418 800
rect 118606 0 118662 800
rect 123850 0 123906 800
rect 129094 0 129150 800
rect 134338 0 134394 800
rect 139582 0 139638 800
rect 144826 0 144882 800
rect 150070 0 150126 800
rect 155314 0 155370 800
rect 160558 0 160614 800
<< obsm2 >>
rect 3240 856 161072 157797
rect 3350 734 8426 856
rect 8594 734 13670 856
rect 13838 734 18914 856
rect 19082 734 24158 856
rect 24326 734 29402 856
rect 29570 734 34646 856
rect 34814 734 39890 856
rect 40058 734 45134 856
rect 45302 734 50378 856
rect 50546 734 55622 856
rect 55790 734 60866 856
rect 61034 734 66110 856
rect 66278 734 71354 856
rect 71522 734 76598 856
rect 76766 734 81842 856
rect 82010 734 87086 856
rect 87254 734 92330 856
rect 92498 734 97574 856
rect 97742 734 102818 856
rect 102986 734 108062 856
rect 108230 734 113306 856
rect 113474 734 118550 856
rect 118718 734 123794 856
rect 123962 734 129038 856
rect 129206 734 134282 856
rect 134450 734 139526 856
rect 139694 734 144770 856
rect 144938 734 150014 856
rect 150182 734 155258 856
rect 155426 734 160502 856
rect 160670 734 161072 856
<< obsm3 >>
rect 4210 2143 158126 157793
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 45875 3435 50208 81837
rect 50688 3435 65568 81837
rect 66048 3435 80928 81837
rect 81408 3435 96288 81837
rect 96768 3435 111648 81837
rect 112128 3435 113837 81837
<< labels >>
rlabel metal2 s 3238 0 3294 800 6 clk
port 1 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 done
port 2 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 reset
port 3 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 serial_line_data[0]
port 4 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 serial_line_data[1]
port 5 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 serial_line_data[2]
port 6 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 serial_line_data[3]
port 7 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 serial_line_data[4]
port 8 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 serial_line_data[5]
port 9 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 serial_line_data[6]
port 10 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 serial_line_data[7]
port 11 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 serial_line_valid
port 12 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 serial_result[0]
port 13 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 serial_result[1]
port 14 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 serial_result[2]
port 15 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 serial_result[3]
port 16 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 serial_result[4]
port 17 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 serial_result[5]
port 18 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 serial_result[6]
port 19 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 serial_result[7]
port 20 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 serial_result_valid
port 21 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 serial_weight_data[0]
port 22 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 serial_weight_data[1]
port 23 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 serial_weight_data[2]
port 24 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 serial_weight_data[3]
port 25 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 serial_weight_data[4]
port 26 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 serial_weight_data[5]
port 27 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 serial_weight_data[6]
port 28 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 serial_weight_data[7]
port 29 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 serial_weight_valid
port 30 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 start
port 31 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 33 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 164000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 23553138
string GDS_FILE /home/kgubbi/kws_final_final/openlane/kws_final_final/runs/24_06_02_21_40/results/signoff/CNN_Accelerator_Top.magic.gds
string GDS_START 1063100
<< end >>


// This is the unpowered netlist.
module CNN_Accelerator_Top (clk,
    done,
    reset,
    serial_line_valid,
    serial_result_valid,
    serial_weight_valid,
    start,
    serial_line_data,
    serial_result,
    serial_weight_data);
 input clk;
 output done;
 input reset;
 input serial_line_valid;
 output serial_result_valid;
 input serial_weight_valid;
 input start;
 input [7:0] serial_line_data;
 output [7:0] serial_result;
 input [7:0] serial_weight_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \control_fsm.line_data[0] ;
 wire \control_fsm.line_data[1] ;
 wire \control_fsm.line_data[2] ;
 wire \control_fsm.line_data[3] ;
 wire \control_fsm.line_data[4] ;
 wire \control_fsm.line_data[5] ;
 wire \control_fsm.line_data[6] ;
 wire \control_fsm.line_data[7] ;
 wire \control_fsm.line_write_addr[0] ;
 wire \control_fsm.line_write_addr[1] ;
 wire \control_fsm.line_write_addr[2] ;
 wire \control_fsm.line_write_addr[3] ;
 wire \control_fsm.line_write_enable ;
 wire \control_fsm.next_state[0] ;
 wire \control_fsm.next_state[1] ;
 wire \control_fsm.next_state[2] ;
 wire \control_fsm.state[0] ;
 wire \control_fsm.state[1] ;
 wire \control_fsm.state[2] ;
 wire \control_fsm.weight_data[0] ;
 wire \control_fsm.weight_data[1] ;
 wire \control_fsm.weight_data[2] ;
 wire \control_fsm.weight_data[3] ;
 wire \control_fsm.weight_data[4] ;
 wire \control_fsm.weight_data[5] ;
 wire \control_fsm.weight_data[6] ;
 wire \control_fsm.weight_data[7] ;
 wire \control_fsm.weight_write_addr[0] ;
 wire \control_fsm.weight_write_addr[1] ;
 wire \control_fsm.weight_write_addr[2] ;
 wire \control_fsm.weight_write_addr[3] ;
 wire \control_fsm.weight_write_enable ;
 wire \line_buffer.data_out[0] ;
 wire \line_buffer.data_out[100] ;
 wire \line_buffer.data_out[101] ;
 wire \line_buffer.data_out[102] ;
 wire \line_buffer.data_out[103] ;
 wire \line_buffer.data_out[104] ;
 wire \line_buffer.data_out[105] ;
 wire \line_buffer.data_out[106] ;
 wire \line_buffer.data_out[107] ;
 wire \line_buffer.data_out[108] ;
 wire \line_buffer.data_out[109] ;
 wire \line_buffer.data_out[10] ;
 wire \line_buffer.data_out[110] ;
 wire \line_buffer.data_out[111] ;
 wire \line_buffer.data_out[112] ;
 wire \line_buffer.data_out[113] ;
 wire \line_buffer.data_out[114] ;
 wire \line_buffer.data_out[115] ;
 wire \line_buffer.data_out[116] ;
 wire \line_buffer.data_out[117] ;
 wire \line_buffer.data_out[118] ;
 wire \line_buffer.data_out[119] ;
 wire \line_buffer.data_out[11] ;
 wire \line_buffer.data_out[120] ;
 wire \line_buffer.data_out[121] ;
 wire \line_buffer.data_out[122] ;
 wire \line_buffer.data_out[123] ;
 wire \line_buffer.data_out[124] ;
 wire \line_buffer.data_out[125] ;
 wire \line_buffer.data_out[126] ;
 wire \line_buffer.data_out[127] ;
 wire \line_buffer.data_out[12] ;
 wire \line_buffer.data_out[13] ;
 wire \line_buffer.data_out[14] ;
 wire \line_buffer.data_out[15] ;
 wire \line_buffer.data_out[16] ;
 wire \line_buffer.data_out[17] ;
 wire \line_buffer.data_out[18] ;
 wire \line_buffer.data_out[19] ;
 wire \line_buffer.data_out[1] ;
 wire \line_buffer.data_out[20] ;
 wire \line_buffer.data_out[21] ;
 wire \line_buffer.data_out[22] ;
 wire \line_buffer.data_out[23] ;
 wire \line_buffer.data_out[24] ;
 wire \line_buffer.data_out[25] ;
 wire \line_buffer.data_out[26] ;
 wire \line_buffer.data_out[27] ;
 wire \line_buffer.data_out[28] ;
 wire \line_buffer.data_out[29] ;
 wire \line_buffer.data_out[2] ;
 wire \line_buffer.data_out[30] ;
 wire \line_buffer.data_out[31] ;
 wire \line_buffer.data_out[32] ;
 wire \line_buffer.data_out[33] ;
 wire \line_buffer.data_out[34] ;
 wire \line_buffer.data_out[35] ;
 wire \line_buffer.data_out[36] ;
 wire \line_buffer.data_out[37] ;
 wire \line_buffer.data_out[38] ;
 wire \line_buffer.data_out[39] ;
 wire \line_buffer.data_out[3] ;
 wire \line_buffer.data_out[40] ;
 wire \line_buffer.data_out[41] ;
 wire \line_buffer.data_out[42] ;
 wire \line_buffer.data_out[43] ;
 wire \line_buffer.data_out[44] ;
 wire \line_buffer.data_out[45] ;
 wire \line_buffer.data_out[46] ;
 wire \line_buffer.data_out[47] ;
 wire \line_buffer.data_out[48] ;
 wire \line_buffer.data_out[49] ;
 wire \line_buffer.data_out[4] ;
 wire \line_buffer.data_out[50] ;
 wire \line_buffer.data_out[51] ;
 wire \line_buffer.data_out[52] ;
 wire \line_buffer.data_out[53] ;
 wire \line_buffer.data_out[54] ;
 wire \line_buffer.data_out[55] ;
 wire \line_buffer.data_out[56] ;
 wire \line_buffer.data_out[57] ;
 wire \line_buffer.data_out[58] ;
 wire \line_buffer.data_out[59] ;
 wire \line_buffer.data_out[5] ;
 wire \line_buffer.data_out[60] ;
 wire \line_buffer.data_out[61] ;
 wire \line_buffer.data_out[62] ;
 wire \line_buffer.data_out[63] ;
 wire \line_buffer.data_out[64] ;
 wire \line_buffer.data_out[65] ;
 wire \line_buffer.data_out[66] ;
 wire \line_buffer.data_out[67] ;
 wire \line_buffer.data_out[68] ;
 wire \line_buffer.data_out[69] ;
 wire \line_buffer.data_out[6] ;
 wire \line_buffer.data_out[70] ;
 wire \line_buffer.data_out[71] ;
 wire \line_buffer.data_out[72] ;
 wire \line_buffer.data_out[73] ;
 wire \line_buffer.data_out[74] ;
 wire \line_buffer.data_out[75] ;
 wire \line_buffer.data_out[76] ;
 wire \line_buffer.data_out[77] ;
 wire \line_buffer.data_out[78] ;
 wire \line_buffer.data_out[79] ;
 wire \line_buffer.data_out[7] ;
 wire \line_buffer.data_out[80] ;
 wire \line_buffer.data_out[81] ;
 wire \line_buffer.data_out[82] ;
 wire \line_buffer.data_out[83] ;
 wire \line_buffer.data_out[84] ;
 wire \line_buffer.data_out[85] ;
 wire \line_buffer.data_out[86] ;
 wire \line_buffer.data_out[87] ;
 wire \line_buffer.data_out[88] ;
 wire \line_buffer.data_out[89] ;
 wire \line_buffer.data_out[8] ;
 wire \line_buffer.data_out[90] ;
 wire \line_buffer.data_out[91] ;
 wire \line_buffer.data_out[92] ;
 wire \line_buffer.data_out[93] ;
 wire \line_buffer.data_out[94] ;
 wire \line_buffer.data_out[95] ;
 wire \line_buffer.data_out[96] ;
 wire \line_buffer.data_out[97] ;
 wire \line_buffer.data_out[98] ;
 wire \line_buffer.data_out[99] ;
 wire \line_buffer.data_out[9] ;
 wire \mac_array.mac[0].mac_unit.b[0] ;
 wire \mac_array.mac[0].mac_unit.b[1] ;
 wire \mac_array.mac[0].mac_unit.b[2] ;
 wire \mac_array.mac[0].mac_unit.b[3] ;
 wire \mac_array.mac[0].mac_unit.b[4] ;
 wire \mac_array.mac[0].mac_unit.b[5] ;
 wire \mac_array.mac[0].mac_unit.b[6] ;
 wire \mac_array.mac[0].mac_unit.b[7] ;
 wire \mac_array.mac[10].mac_unit.b[0] ;
 wire \mac_array.mac[10].mac_unit.b[1] ;
 wire \mac_array.mac[10].mac_unit.b[2] ;
 wire \mac_array.mac[10].mac_unit.b[3] ;
 wire \mac_array.mac[10].mac_unit.b[4] ;
 wire \mac_array.mac[10].mac_unit.b[5] ;
 wire \mac_array.mac[10].mac_unit.b[6] ;
 wire \mac_array.mac[10].mac_unit.b[7] ;
 wire \mac_array.mac[11].mac_unit.b[0] ;
 wire \mac_array.mac[11].mac_unit.b[1] ;
 wire \mac_array.mac[11].mac_unit.b[2] ;
 wire \mac_array.mac[11].mac_unit.b[3] ;
 wire \mac_array.mac[11].mac_unit.b[4] ;
 wire \mac_array.mac[11].mac_unit.b[5] ;
 wire \mac_array.mac[11].mac_unit.b[6] ;
 wire \mac_array.mac[11].mac_unit.b[7] ;
 wire \mac_array.mac[12].mac_unit.b[0] ;
 wire \mac_array.mac[12].mac_unit.b[1] ;
 wire \mac_array.mac[12].mac_unit.b[2] ;
 wire \mac_array.mac[12].mac_unit.b[3] ;
 wire \mac_array.mac[12].mac_unit.b[4] ;
 wire \mac_array.mac[12].mac_unit.b[5] ;
 wire \mac_array.mac[12].mac_unit.b[6] ;
 wire \mac_array.mac[12].mac_unit.b[7] ;
 wire \mac_array.mac[13].mac_unit.b[0] ;
 wire \mac_array.mac[13].mac_unit.b[1] ;
 wire \mac_array.mac[13].mac_unit.b[2] ;
 wire \mac_array.mac[13].mac_unit.b[3] ;
 wire \mac_array.mac[13].mac_unit.b[4] ;
 wire \mac_array.mac[13].mac_unit.b[5] ;
 wire \mac_array.mac[13].mac_unit.b[6] ;
 wire \mac_array.mac[13].mac_unit.b[7] ;
 wire \mac_array.mac[14].mac_unit.b[0] ;
 wire \mac_array.mac[14].mac_unit.b[1] ;
 wire \mac_array.mac[14].mac_unit.b[2] ;
 wire \mac_array.mac[14].mac_unit.b[3] ;
 wire \mac_array.mac[14].mac_unit.b[4] ;
 wire \mac_array.mac[14].mac_unit.b[5] ;
 wire \mac_array.mac[14].mac_unit.b[6] ;
 wire \mac_array.mac[14].mac_unit.b[7] ;
 wire \mac_array.mac[15].mac_unit.b[0] ;
 wire \mac_array.mac[15].mac_unit.b[1] ;
 wire \mac_array.mac[15].mac_unit.b[2] ;
 wire \mac_array.mac[15].mac_unit.b[3] ;
 wire \mac_array.mac[15].mac_unit.b[4] ;
 wire \mac_array.mac[15].mac_unit.b[5] ;
 wire \mac_array.mac[15].mac_unit.b[6] ;
 wire \mac_array.mac[15].mac_unit.b[7] ;
 wire \mac_array.mac[1].mac_unit.b[0] ;
 wire \mac_array.mac[1].mac_unit.b[1] ;
 wire \mac_array.mac[1].mac_unit.b[2] ;
 wire \mac_array.mac[1].mac_unit.b[3] ;
 wire \mac_array.mac[1].mac_unit.b[4] ;
 wire \mac_array.mac[1].mac_unit.b[5] ;
 wire \mac_array.mac[1].mac_unit.b[6] ;
 wire \mac_array.mac[1].mac_unit.b[7] ;
 wire \mac_array.mac[2].mac_unit.b[0] ;
 wire \mac_array.mac[2].mac_unit.b[1] ;
 wire \mac_array.mac[2].mac_unit.b[2] ;
 wire \mac_array.mac[2].mac_unit.b[3] ;
 wire \mac_array.mac[2].mac_unit.b[4] ;
 wire \mac_array.mac[2].mac_unit.b[5] ;
 wire \mac_array.mac[2].mac_unit.b[6] ;
 wire \mac_array.mac[2].mac_unit.b[7] ;
 wire \mac_array.mac[3].mac_unit.b[0] ;
 wire \mac_array.mac[3].mac_unit.b[1] ;
 wire \mac_array.mac[3].mac_unit.b[2] ;
 wire \mac_array.mac[3].mac_unit.b[3] ;
 wire \mac_array.mac[3].mac_unit.b[4] ;
 wire \mac_array.mac[3].mac_unit.b[5] ;
 wire \mac_array.mac[3].mac_unit.b[6] ;
 wire \mac_array.mac[3].mac_unit.b[7] ;
 wire \mac_array.mac[4].mac_unit.b[0] ;
 wire \mac_array.mac[4].mac_unit.b[1] ;
 wire \mac_array.mac[4].mac_unit.b[2] ;
 wire \mac_array.mac[4].mac_unit.b[3] ;
 wire \mac_array.mac[4].mac_unit.b[4] ;
 wire \mac_array.mac[4].mac_unit.b[5] ;
 wire \mac_array.mac[4].mac_unit.b[6] ;
 wire \mac_array.mac[4].mac_unit.b[7] ;
 wire \mac_array.mac[5].mac_unit.b[0] ;
 wire \mac_array.mac[5].mac_unit.b[1] ;
 wire \mac_array.mac[5].mac_unit.b[2] ;
 wire \mac_array.mac[5].mac_unit.b[3] ;
 wire \mac_array.mac[5].mac_unit.b[4] ;
 wire \mac_array.mac[5].mac_unit.b[5] ;
 wire \mac_array.mac[5].mac_unit.b[6] ;
 wire \mac_array.mac[5].mac_unit.b[7] ;
 wire \mac_array.mac[6].mac_unit.b[0] ;
 wire \mac_array.mac[6].mac_unit.b[1] ;
 wire \mac_array.mac[6].mac_unit.b[2] ;
 wire \mac_array.mac[6].mac_unit.b[3] ;
 wire \mac_array.mac[6].mac_unit.b[4] ;
 wire \mac_array.mac[6].mac_unit.b[5] ;
 wire \mac_array.mac[6].mac_unit.b[6] ;
 wire \mac_array.mac[6].mac_unit.b[7] ;
 wire \mac_array.mac[7].mac_unit.b[0] ;
 wire \mac_array.mac[7].mac_unit.b[1] ;
 wire \mac_array.mac[7].mac_unit.b[2] ;
 wire \mac_array.mac[7].mac_unit.b[3] ;
 wire \mac_array.mac[7].mac_unit.b[4] ;
 wire \mac_array.mac[7].mac_unit.b[5] ;
 wire \mac_array.mac[7].mac_unit.b[6] ;
 wire \mac_array.mac[7].mac_unit.b[7] ;
 wire \mac_array.mac[8].mac_unit.b[0] ;
 wire \mac_array.mac[8].mac_unit.b[1] ;
 wire \mac_array.mac[8].mac_unit.b[2] ;
 wire \mac_array.mac[8].mac_unit.b[3] ;
 wire \mac_array.mac[8].mac_unit.b[4] ;
 wire \mac_array.mac[8].mac_unit.b[5] ;
 wire \mac_array.mac[8].mac_unit.b[6] ;
 wire \mac_array.mac[8].mac_unit.b[7] ;
 wire \mac_array.mac[9].mac_unit.b[0] ;
 wire \mac_array.mac[9].mac_unit.b[1] ;
 wire \mac_array.mac[9].mac_unit.b[2] ;
 wire \mac_array.mac[9].mac_unit.b[3] ;
 wire \mac_array.mac[9].mac_unit.b[4] ;
 wire \mac_array.mac[9].mac_unit.b[5] ;
 wire \mac_array.mac[9].mac_unit.b[6] ;
 wire \mac_array.mac[9].mac_unit.b[7] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net242;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net243;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net244;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net245;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net246;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net247;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net248;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net249;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net25;
 wire net250;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net251;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net252;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net253;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net254;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net255;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net256;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net257;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net258;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net259;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net26;
 wire net260;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net261;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net262;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net263;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net264;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net265;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net266;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net267;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net268;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net269;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net27;
 wire net270;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net271;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net272;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net273;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net274;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net275;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net276;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net277;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2777;
 wire net2779;
 wire net278;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net279;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net28;
 wire net280;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net281;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net282;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net283;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net284;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net285;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net286;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net287;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net288;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net289;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net29;
 wire net290;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net291;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net292;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net293;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net294;
 wire net2940;
 wire net2941;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net295;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net296;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net297;
 wire net2970;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net298;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net299;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3;
 wire net30;
 wire net300;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net301;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net302;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net303;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net304;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net305;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net306;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net307;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net308;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net309;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net31;
 wire net310;
 wire net3100;
 wire net3101;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net311;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net312;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net313;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net314;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net315;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net316;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net317;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net318;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net319;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net32;
 wire net320;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net321;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3214;
 wire net3215;
 wire net3219;
 wire net322;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net323;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net324;
 wire net3240;
 wire net3241;
 wire net3243;
 wire net3244;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net325;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net326;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net327;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net328;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net329;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net33;
 wire net330;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net331;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net332;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net333;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net334;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net335;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net336;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net337;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net338;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net339;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net34;
 wire net340;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net341;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net342;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net343;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net344;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net345;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net346;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net347;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net348;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net349;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net35;
 wire net350;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net351;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net352;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net353;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net354;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net355;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3558;
 wire net3559;
 wire net356;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3569;
 wire net357;
 wire net3570;
 wire net3571;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net358;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net359;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net36;
 wire net360;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net361;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net362;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net363;
 wire net3630;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net364;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net365;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net366;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net367;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net368;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net369;
 wire net3690;
 wire net3694;
 wire net3695;
 wire net3698;
 wire net3699;
 wire net37;
 wire net370;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net371;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3716;
 wire net3719;
 wire net372;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net373;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net374;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net375;
 wire net3750;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net376;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3769;
 wire net377;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net378;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net379;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net38;
 wire net380;
 wire net3809;
 wire net381;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net382;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net383;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net384;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net385;
 wire net3851;
 wire net3858;
 wire net3859;
 wire net386;
 wire net3860;
 wire net3861;
 wire net3868;
 wire net3869;
 wire net387;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net388;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \next_state[0] ;
 wire \result[0][0] ;
 wire \result[0][1] ;
 wire \result[0][2] ;
 wire \result[0][3] ;
 wire \result[0][4] ;
 wire \result[0][5] ;
 wire \result[0][6] ;
 wire \result[0][7] ;
 wire \result[10][0] ;
 wire \result[10][1] ;
 wire \result[10][2] ;
 wire \result[10][3] ;
 wire \result[10][4] ;
 wire \result[10][5] ;
 wire \result[10][6] ;
 wire \result[10][7] ;
 wire \result[11][0] ;
 wire \result[11][1] ;
 wire \result[11][2] ;
 wire \result[11][3] ;
 wire \result[11][4] ;
 wire \result[11][5] ;
 wire \result[11][6] ;
 wire \result[11][7] ;
 wire \result[13][0] ;
 wire \result[13][1] ;
 wire \result[13][2] ;
 wire \result[13][3] ;
 wire \result[13][4] ;
 wire \result[13][5] ;
 wire \result[13][6] ;
 wire \result[13][7] ;
 wire \result_index[0] ;
 wire \result_index[1] ;
 wire \result_index[2] ;
 wire \result_index[3] ;
 wire \state[0] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_06462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__06478__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__C (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A1 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A0 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__A0 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__A0 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06495__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06495__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06496__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06496__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06497__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06497__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__A1 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06501__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06501__S (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__C_N (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06506__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06506__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__S (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__A (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06515__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A0 (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A1 (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__06518__A0 (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__06519__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06520__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06520__A1 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__A_N (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A_N (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__A1 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06528__A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06530__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__A1 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06538__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06538__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__S (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06549__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06549__S (.DIODE(_00681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06554__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06554__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__S (.DIODE(_00682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__B (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A_N (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__A1 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__A0 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__A0 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__A0 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__S (.DIODE(_00684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06570__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06570__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06571__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06571__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06573__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06573__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__S (.DIODE(_00685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06578__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A1 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A1 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__S (.DIODE(_00686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A1 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__A_N (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A0 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A1 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__A1 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A1 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__S (.DIODE(_00689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A1 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__A (.DIODE(_00674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__S (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__A_N (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__B (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__A_N (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__B (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__A1 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__A1 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__B2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__B (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__B2 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__C (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__B2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A1_N (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06711__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__B2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__C (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A1_N (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A1 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__B2 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A1 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A1 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B2 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__B2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__A1 (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__B2 (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__B (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__B2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B2 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__B (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__B (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__B2 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__B (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__C (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A1_N (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__B (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__B2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__B2 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__B2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__B2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A1 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__B2 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__B2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__B (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B2 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__B (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B2 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__D (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__B2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A1 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A2 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__B (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__D (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A1 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B2 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__B (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A2 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A1 (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__D (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A1 (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__D (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__B1 (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__B2 (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__B1 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__D (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B1 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__C (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__D (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A2 (.DIODE(net2066));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__D (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A1 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__C (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A1_N (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__B (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A1 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B2 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__B2 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__B2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A1 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A1 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__B2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A1 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B2 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__B (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B2 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B2 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A1 (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__B (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A1 (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__B2 (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__A1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__B2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__B (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A1 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A2 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__B (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A1 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B2 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B2 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A2 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__B2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A1 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A2 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A1 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A2 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__B (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A1 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A2 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__D (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A1 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__B1 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__B2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__D (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A2_N (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B2 (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A1 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B2 (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__B1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__D (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A2 (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__B2 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__B (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__D (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__A2 (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__D (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A1 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__B (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A2 (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__B (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A2 (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A1 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__B (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__B (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__C (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07867__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A1 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A2 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B2 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__B (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__D (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B2 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__B (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A1 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__B (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A1 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__B1 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__B (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__B2 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A (.DIODE(_02075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A1 (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A1 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B2 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__B2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A1 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__B2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__A1 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__B2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__B (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B2 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__B (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__C (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A1_N (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__D (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B1 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__C (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A1 (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__B (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A2 (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__B2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A1 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__B2 (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__B (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A1 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B2 (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__C (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A1_N (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__B2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B2 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__B (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A1 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__D (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A2 (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__D (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A2_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A2 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08516__A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__C (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B1 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A1 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__C (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__C (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A1_N (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__08569__B (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A2 (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__B1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__C (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__D (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A1_N (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A2_N (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__A1 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__B2 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08622__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__B (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A1 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__B (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__C (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__C1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__B (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__B (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A2 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__B (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__C (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__A1 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__B (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__B (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A1 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B2 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__B (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A1 (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A2 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__C (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__C (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__B2 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__C (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__D (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__B1 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__C (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__D (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__B1 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__C (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__D (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A1 (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__C (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A2 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B1 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1_N (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__A2 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__B1 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__C (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__D (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__B (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__B (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__C (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A1 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A2 (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B (.DIODE(_02973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__C (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08912__A (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__A1 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__A2 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08913__B1 (.DIODE(_02973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__B (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__B1 (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__B (.DIODE(_02996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__B (.DIODE(_03019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A2 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__B1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__C (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__B (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(_03061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__B (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A1 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A2 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A2 (.DIODE(_03108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__B1 (.DIODE(_03100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__B (.DIODE(_03108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B (.DIODE(_03137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__B (.DIODE(_03137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__B (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__B (.DIODE(_03144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A (.DIODE(_03192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__B (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A1 (.DIODE(_02087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A_N (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__B (.DIODE(_03205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A (.DIODE(_03210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__A1 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__09177__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A0 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A0 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__A0 (.DIODE(net2286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__09183__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09189__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A0 (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A0 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A0 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__S (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A0 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A0 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__S (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__S (.DIODE(_03246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A1 (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A1 (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__S (.DIODE(_03248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09248__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__S (.DIODE(_03250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__S (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A0 (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__S (.DIODE(_03254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A1 (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A0 (.DIODE(net1681));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A0 (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09292__S (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A1 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__S (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__A1 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A1 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A1 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__A1 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A1 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A1 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A1 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__S (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__A0 (.DIODE(net2367));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A0 (.DIODE(net1874));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__A0 (.DIODE(net2326));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A0 (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A0 (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA__09320__A0 (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A1 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A1 (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__S (.DIODE(_03262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__B1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B1 (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__B1 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__S (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__B (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__C (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A2 (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B (.DIODE(_03265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A0 (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A0 (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A0 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A0 (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A0 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__S (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__C (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__B1 (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A2 (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__B (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__C (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__B (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A1 (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__D (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A2_N (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B2 (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__A2 (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B2 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__B (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A2 (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__D (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B2 (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A1 (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B1 (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A1 (.DIODE(net2511));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__B2 (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__C (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A1_N (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A2 (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09638__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09654__B2 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__B2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__B (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__B (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__C (.DIODE(net2459));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__A2 (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__B (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__A1 (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__A2 (.DIODE(net2459));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__B2 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__B (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__C (.DIODE(net2459));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A2 (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A2 (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__B2 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__B2 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__C (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A1_N (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A2_N (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A2 (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__B (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A1 (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__D (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__A (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__A1 (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__B1 (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__B2 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__B (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09852__A1 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__C (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__D (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A1_N (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A2_N (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__B (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__B (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__B (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__C (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__C (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__A2 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10022__A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A2 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__D (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__D (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__D (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__B (.DIODE(_03780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__B (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A1 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__B2 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A1 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__B2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A1 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__B2 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__B2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__B2 (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10399__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__B1 (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__D (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__D (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__B1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__C (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__B (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__B2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A2 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A1 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A1 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__B (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__B2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A4 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__A1 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__A2 (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__B (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__C (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A1 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A2 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A1 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B2 (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A1 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__B2 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__B (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A2 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A1 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__B2 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__B (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__C (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__D (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A1 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A2 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__C1 (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__A2 (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__B (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B1 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B2 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__C (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A1 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A1 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A2 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__B2 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__B (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A2 (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B1 (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B2 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__A1 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__B1 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__B2 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__D (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__B (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A1 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__B2 (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A1 (.DIODE(_04568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A2 (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__C (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A2 (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A2 (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__C (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__C (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__D (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__B1 (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__D (.DIODE(net675));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__A1 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__A2 (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__B1 (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__B2 (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A1 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A2 (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A3 (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A4 (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__B (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__A2 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__B (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__B (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A2 (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__B (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__C (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__C (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__C (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__C (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__B (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__B2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__B1 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__D (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__D (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__B (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A2 (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__B (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__C (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__B (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A1 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A2 (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__B (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__10842__C (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10842__D (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1_N (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A2_N (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A2 (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__A2 (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__B (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__B (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A1 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__B (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A2 (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__B (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__B2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__C (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A1_N (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A1 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__C1 (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__A2 (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A2 (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A1 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__B2 (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A1 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A2 (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A1 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__B (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__B2 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__B (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__A2 (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__B2 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__C (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__A2 (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__A (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A1 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__B (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A1 (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__B2 (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__B2 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__B2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__A1 (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__B (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__B (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__B (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__B2 (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__B (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__B (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__B2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__D (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__C (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A1_N (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__B (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__B1 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A1 (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__C (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A1 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A2 (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__B2 (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__C (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1_N (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A1 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11341__B (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__C (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A1_N (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__B1 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A1 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__B (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__B2 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__B (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A1 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A2 (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A2 (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__B2 (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__B (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A1 (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A1_N (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__A2 (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A2 (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__A (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__A2 (.DIODE(_05500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A (.DIODE(_04568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__B (.DIODE(_05560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11667__A (.DIODE(_05567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__A (.DIODE(_05581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A (.DIODE(_05581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A (.DIODE(_05581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__B1 (.DIODE(_05560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__A (.DIODE(_05611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__A (.DIODE(_05622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__A1 (.DIODE(_05622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B (.DIODE(_05642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__A2 (.DIODE(_05642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__B (.DIODE(_05729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__B (.DIODE(_05733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__B (.DIODE(_05745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__B1 (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__B2 (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A2 (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__B (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B (.DIODE(_05837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A1 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A2 (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__B2 (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__B (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__B2 (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__C (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__B2 (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__B1 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__12130__A1_N (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A2 (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__C (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B2 (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__A (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__C (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A2 (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A2 (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A1 (.DIODE(_06255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__B2 (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A1 (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__B1 (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A1 (.DIODE(_06300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12429__A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A1 (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__C (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__D (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__B1 (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__B2 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A1_N (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__A2_N (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__B (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__B2 (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__D (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12475__A2_N (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12477__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12481__B2 (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__B2 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__C (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A2 (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__A (.DIODE(_03518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A2 (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__C1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__B (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__B (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__B (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__C (.DIODE(net2635));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__A (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__B (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__B2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__B (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__B (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__B2 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A0 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__S (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__B1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__B1 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__B1 (.DIODE(_06448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12579__B1 (.DIODE(_06451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__B1 (.DIODE(net2635));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__B1 (.DIODE(_06454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__B1 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__A1 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12589__B1 (.DIODE(net2635));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__B1 (.DIODE(net2635));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A_N (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__B (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__B1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A1 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A1 (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__A3 (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__S0 (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__S1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__A1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__S (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A0 (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__A0 (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A0 (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__A0 (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__12603__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__A0 (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A0 (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A0 (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__A0 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__S (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12608__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12624__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12626__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12632__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12651__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12653__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12682__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12721__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12737__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12747__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12749__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12763__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12765__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12777__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12789__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12872__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12891__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12893__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12895__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12909__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12913__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12915__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12920__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12925__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12929__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12931__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12932__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12933__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12935__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12937__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12939__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12943__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__CLK (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__CLK (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net2459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net2066));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net2367));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net1874));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net2326));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net1681));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net2286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(net2511));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1037_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1251_A (.DIODE(_00673_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1278_A (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1317_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1323_A (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1350_A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1472_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1547_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1582_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1587_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1665_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1712_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1823_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1846_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1858_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1896_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1909_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1918_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1928_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1960_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1974_A (.DIODE(net941));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1985_A (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2005_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2048_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2058_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2077_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2083_A (.DIODE(net800));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2117_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2147_A (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2211_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2223_A (.DIODE(net767));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2228_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2239_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2261_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2285_A (.DIODE(net899));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2291_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2303_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2326_A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2368_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2374_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2396_A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2401_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2417_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2430_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2435_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2440_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2448_A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2491_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2497_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2503_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2509_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2638_A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2666_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2762_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2785_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2946_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3016_A (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3020_A (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3033_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3103_A (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3181_A (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3211_A (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3216_A (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3224_A (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3232_A (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3282_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3297_A (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3339_A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3343_A (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3353_A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3369_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3371_A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3381_A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3409_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3419_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3425_A (.DIODE(net797));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3509_A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3546_A (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3587_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold814_A (.DIODE(_03267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_202_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_208_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_212_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_214_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_214_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_218_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_220_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_222_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_224_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_224_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_226_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_230_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_230_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_232_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_234_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_236_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_236_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_238_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_240_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_240_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_244_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_244_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_246_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_246_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_248_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_248_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_250_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_252_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_252_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_254_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_254_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_256_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_258_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_260_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_260_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_262_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_264_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_264_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_266_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_268_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_270_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_270_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_271_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_272_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_272_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_274_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_274_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_276_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_276_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_277_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_278_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_279_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_280_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_280_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_282_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_282_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_284_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_284_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_285_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_285_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_285_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_285_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06476_ (.A(net714),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_2 _06477_ (.A(net19),
    .Y(_00666_));
 sky130_fd_sc_hd__inv_2 _06478_ (.A(net10),
    .Y(_00667_));
 sky130_fd_sc_hd__inv_2 _06479_ (.A(net1114),
    .Y(_00668_));
 sky130_fd_sc_hd__inv_2 _06480_ (.A(net1021),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_2 _06481_ (.A(net203),
    .Y(_00000_));
 sky130_fd_sc_hd__or3b_1 _06482_ (.A(net1192),
    .B(net1401),
    .C_N(net1337),
    .X(_00670_));
 sky130_fd_sc_hd__nor3_1 _06483_ (.A(net1621),
    .B(net1460),
    .C(net1402),
    .Y(_00671_));
 sky130_fd_sc_hd__mux2_1 _06484_ (.A0(net1448),
    .A1(net174),
    .S(net33),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _06485_ (.A0(net1488),
    .A1(net175),
    .S(net33),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _06486_ (.A0(net2495),
    .A1(net2287),
    .S(net33),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _06487_ (.A0(net2489),
    .A1(net1014),
    .S(net33),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _06488_ (.A0(net1861),
    .A1(net1018),
    .S(net33),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(net1686),
    .A1(net179),
    .S(net33),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _06490_ (.A0(net1652),
    .A1(net180),
    .S(net33),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _06491_ (.A0(net1574),
    .A1(net181),
    .S(net33),
    .X(_00657_));
 sky130_fd_sc_hd__and3b_4 _06492_ (.A_N(net1520),
    .B(net1444),
    .C(net1337),
    .X(_00672_));
 sky130_fd_sc_hd__or3b_2 _06493_ (.A(net1433),
    .B(net1460),
    .C_N(_00672_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _06494_ (.A0(net174),
    .A1(net1429),
    .S(net1461),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _06495_ (.A0(net175),
    .A1(net473),
    .S(net1461),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _06496_ (.A0(net2287),
    .A1(net2455),
    .S(net1461),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _06497_ (.A0(net1014),
    .A1(net2101),
    .S(net1461),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _06498_ (.A0(net1018),
    .A1(net1825),
    .S(net1461),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _06499_ (.A0(net179),
    .A1(net2961),
    .S(net1461),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _06500_ (.A0(net180),
    .A1(net914),
    .S(net1461),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _06501_ (.A0(net181),
    .A1(net731),
    .S(net1461),
    .X(_00649_));
 sky130_fd_sc_hd__and3b_4 _06502_ (.A_N(net1444),
    .B(net1520),
    .C(net1337),
    .X(_00674_));
 sky130_fd_sc_hd__or3b_1 _06503_ (.A(net1433),
    .B(net1460),
    .C_N(_00674_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _06504_ (.A0(net174),
    .A1(net1393),
    .S(net1434),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _06505_ (.A0(net175),
    .A1(net440),
    .S(net1434),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _06506_ (.A0(net2287),
    .A1(net2385),
    .S(net1434),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _06507_ (.A0(net1014),
    .A1(net2262),
    .S(net1434),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _06508_ (.A0(net1018),
    .A1(net1879),
    .S(net1434),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _06509_ (.A0(net179),
    .A1(net1966),
    .S(net1434),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _06510_ (.A0(net180),
    .A1(net1773),
    .S(net1434),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _06511_ (.A0(net181),
    .A1(net1632),
    .S(net1434),
    .X(_00641_));
 sky130_fd_sc_hd__and3_4 _06512_ (.A(net1337),
    .B(net1520),
    .C(net1444),
    .X(_00676_));
 sky130_fd_sc_hd__or3b_4 _06513_ (.A(net1621),
    .B(net1460),
    .C_N(_00676_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _06514_ (.A0(net174),
    .A1(net1425),
    .S(_00677_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _06515_ (.A0(net175),
    .A1(net3043),
    .S(_00677_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _06516_ (.A0(net2287),
    .A1(net2421),
    .S(_00677_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _06517_ (.A0(net1013),
    .A1(net2690),
    .S(_00677_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _06518_ (.A0(net1017),
    .A1(net2848),
    .S(_00677_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _06519_ (.A0(net179),
    .A1(net3432),
    .S(_00677_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _06520_ (.A0(net180),
    .A1(net1752),
    .S(_00677_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _06521_ (.A0(net181),
    .A1(net3230),
    .S(_00677_),
    .X(_00633_));
 sky130_fd_sc_hd__and2b_2 _06522_ (.A_N(net1621),
    .B(net1460),
    .X(_00678_));
 sky130_fd_sc_hd__and2b_1 _06523_ (.A_N(net1402),
    .B(_00678_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _06524_ (.A0(net3628),
    .A1(net174),
    .S(net1403),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _06525_ (.A0(net421),
    .A1(net175),
    .S(net1403),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _06526_ (.A0(net2513),
    .A1(net2287),
    .S(net1403),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _06527_ (.A0(net3563),
    .A1(net1014),
    .S(net1403),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _06528_ (.A0(net2518),
    .A1(net1018),
    .S(net1403),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _06529_ (.A0(net1909),
    .A1(net179),
    .S(net1403),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _06530_ (.A0(net2303),
    .A1(net180),
    .S(net1403),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _06531_ (.A0(net3226),
    .A1(net181),
    .S(net1403),
    .X(_00625_));
 sky130_fd_sc_hd__nand2_4 _06532_ (.A(_00672_),
    .B(_00678_),
    .Y(_00680_));
 sky130_fd_sc_hd__mux2_1 _06533_ (.A0(net174),
    .A1(net1421),
    .S(_00680_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _06534_ (.A0(net175),
    .A1(net1471),
    .S(_00680_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _06535_ (.A0(net2287),
    .A1(net2670),
    .S(_00680_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _06536_ (.A0(net1014),
    .A1(net1995),
    .S(_00680_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _06537_ (.A0(net1018),
    .A1(net2243),
    .S(_00680_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _06538_ (.A0(net179),
    .A1(net1813),
    .S(_00680_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _06539_ (.A0(net180),
    .A1(net1721),
    .S(_00680_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _06540_ (.A0(net181),
    .A1(net1611),
    .S(_00680_),
    .X(_00617_));
 sky130_fd_sc_hd__nand2_4 _06541_ (.A(_00674_),
    .B(_00678_),
    .Y(_00681_));
 sky130_fd_sc_hd__mux2_1 _06542_ (.A0(net174),
    .A1(net1407),
    .S(_00681_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _06543_ (.A0(net175),
    .A1(net1510),
    .S(_00681_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _06544_ (.A0(net2287),
    .A1(net3591),
    .S(_00681_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _06545_ (.A0(net1014),
    .A1(net2438),
    .S(_00681_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _06546_ (.A0(net1018),
    .A1(net2443),
    .S(_00681_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _06547_ (.A0(net179),
    .A1(net3586),
    .S(_00681_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _06548_ (.A0(net180),
    .A1(net3576),
    .S(_00681_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _06549_ (.A0(net181),
    .A1(net3243),
    .S(_00681_),
    .X(_00609_));
 sky130_fd_sc_hd__nand2_4 _06550_ (.A(_00676_),
    .B(_00678_),
    .Y(_00682_));
 sky130_fd_sc_hd__mux2_1 _06551_ (.A0(net174),
    .A1(net3126),
    .S(_00682_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _06552_ (.A0(net175),
    .A1(net3152),
    .S(_00682_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _06553_ (.A0(net2287),
    .A1(net3635),
    .S(_00682_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _06554_ (.A0(net1014),
    .A1(net3629),
    .S(_00682_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _06555_ (.A0(net1018),
    .A1(net3060),
    .S(_00682_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _06556_ (.A0(net179),
    .A1(net3546),
    .S(_00682_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _06557_ (.A0(net180),
    .A1(net3549),
    .S(_00682_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _06558_ (.A0(net181),
    .A1(net3238),
    .S(_00682_),
    .X(_00601_));
 sky130_fd_sc_hd__and2b_4 _06559_ (.A_N(net1460),
    .B(net1621),
    .X(_00683_));
 sky130_fd_sc_hd__and2b_4 _06560_ (.A_N(net1402),
    .B(_00683_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _06561_ (.A0(net1492),
    .A1(net174),
    .S(_00684_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _06562_ (.A0(net1541),
    .A1(net175),
    .S(_00684_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _06563_ (.A0(net1763),
    .A1(net2287),
    .S(_00684_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _06564_ (.A0(net1664),
    .A1(net1014),
    .S(_00684_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _06565_ (.A0(net2311),
    .A1(net1018),
    .S(_00684_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _06566_ (.A0(net1960),
    .A1(net179),
    .S(_00684_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _06567_ (.A0(net1946),
    .A1(net180),
    .S(_00684_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _06568_ (.A0(net1636),
    .A1(net181),
    .S(_00684_),
    .X(_00593_));
 sky130_fd_sc_hd__nand2_4 _06569_ (.A(_00672_),
    .B(_00683_),
    .Y(_00685_));
 sky130_fd_sc_hd__mux2_1 _06570_ (.A0(net174),
    .A1(net1411),
    .S(_00685_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _06571_ (.A0(net175),
    .A1(net1467),
    .S(_00685_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _06572_ (.A0(net2287),
    .A1(net3698),
    .S(_00685_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _06573_ (.A0(net1014),
    .A1(net3719),
    .S(_00685_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _06574_ (.A0(net1018),
    .A1(net3756),
    .S(_00685_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _06575_ (.A0(net179),
    .A1(net3769),
    .S(_00685_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _06576_ (.A0(net180),
    .A1(net1658),
    .S(_00685_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _06577_ (.A0(net181),
    .A1(net1586),
    .S(_00685_),
    .X(_00585_));
 sky130_fd_sc_hd__nand2_4 _06578_ (.A(_00674_),
    .B(_00683_),
    .Y(_00686_));
 sky130_fd_sc_hd__mux2_1 _06579_ (.A0(net174),
    .A1(net1504),
    .S(_00686_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _06580_ (.A0(net175),
    .A1(net1560),
    .S(_00686_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _06581_ (.A0(net2287),
    .A1(net2471),
    .S(_00686_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _06582_ (.A0(net1014),
    .A1(net2272),
    .S(_00686_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _06583_ (.A0(net1018),
    .A1(net2110),
    .S(_00686_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _06584_ (.A0(net179),
    .A1(net2215),
    .S(_00686_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _06585_ (.A0(net180),
    .A1(net2062),
    .S(_00686_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _06586_ (.A0(net181),
    .A1(net3002),
    .S(_00686_),
    .X(_00577_));
 sky130_fd_sc_hd__nand2_4 _06587_ (.A(_00676_),
    .B(_00683_),
    .Y(_00687_));
 sky130_fd_sc_hd__mux2_1 _06588_ (.A0(net174),
    .A1(net1456),
    .S(_00687_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _06589_ (.A0(net175),
    .A1(net1527),
    .S(_00687_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _06590_ (.A0(net2287),
    .A1(net776),
    .S(_00687_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _06591_ (.A0(net1014),
    .A1(net2268),
    .S(_00687_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _06592_ (.A0(net1018),
    .A1(net2293),
    .S(_00687_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _06593_ (.A0(net179),
    .A1(net2170),
    .S(_00687_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _06594_ (.A0(net180),
    .A1(net2138),
    .S(_00687_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _06595_ (.A0(net181),
    .A1(net2943),
    .S(_00687_),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _06596_ (.A(net1621),
    .B(net1460),
    .X(_00688_));
 sky130_fd_sc_hd__and2b_4 _06597_ (.A_N(net1402),
    .B(net1622),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _06598_ (.A0(net1496),
    .A1(net174),
    .S(_00689_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _06599_ (.A0(net1550),
    .A1(net175),
    .S(_00689_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _06600_ (.A0(net2584),
    .A1(net2287),
    .S(_00689_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _06601_ (.A0(net2578),
    .A1(net1014),
    .S(_00689_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _06602_ (.A0(net2590),
    .A1(net1018),
    .S(_00689_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _06603_ (.A0(net2205),
    .A1(net179),
    .S(_00689_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _06604_ (.A0(net2056),
    .A1(net180),
    .S(_00689_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _06605_ (.A0(net1644),
    .A1(net181),
    .S(_00689_),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_4 _06606_ (.A(_00672_),
    .B(net1622),
    .Y(_00690_));
 sky130_fd_sc_hd__mux2_1 _06607_ (.A0(net174),
    .A1(net1385),
    .S(_00690_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _06608_ (.A0(net175),
    .A1(net1482),
    .S(_00690_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _06609_ (.A0(net2287),
    .A1(net1160),
    .S(_00690_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _06610_ (.A0(net1014),
    .A1(net2247),
    .S(_00690_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _06611_ (.A0(net1018),
    .A1(net2258),
    .S(_00690_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _06612_ (.A0(net179),
    .A1(net1792),
    .S(_00690_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _06613_ (.A0(net180),
    .A1(net1757),
    .S(_00690_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _06614_ (.A0(net181),
    .A1(net1603),
    .S(_00690_),
    .X(_00553_));
 sky130_fd_sc_hd__nand2_4 _06615_ (.A(_00674_),
    .B(net1622),
    .Y(_00691_));
 sky130_fd_sc_hd__mux2_1 _06616_ (.A0(net174),
    .A1(net1500),
    .S(_00691_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _06617_ (.A0(net175),
    .A1(net1514),
    .S(_00691_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _06618_ (.A0(net2287),
    .A1(net3581),
    .S(_00691_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _06619_ (.A0(net1014),
    .A1(net3569),
    .S(_00691_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _06620_ (.A0(net1018),
    .A1(net2401),
    .S(_00691_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _06621_ (.A0(net179),
    .A1(net2185),
    .S(_00691_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _06622_ (.A0(net180),
    .A1(net3365),
    .S(_00691_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _06623_ (.A0(net181),
    .A1(net3247),
    .S(_00691_),
    .X(_00545_));
 sky130_fd_sc_hd__and2b_1 _06624_ (.A_N(net1110),
    .B(net1245),
    .X(_00692_));
 sky130_fd_sc_hd__nand2b_1 _06625_ (.A_N(net1110),
    .B(net1245),
    .Y(_00693_));
 sky130_fd_sc_hd__and4_1 _06626_ (.A(net857),
    .B(net938),
    .C(net848),
    .D(net770),
    .X(_00694_));
 sky130_fd_sc_hd__and2_1 _06627_ (.A(net1550),
    .B(net770),
    .X(_00695_));
 sky130_fd_sc_hd__a21oi_1 _06628_ (.A1(net857),
    .A2(net848),
    .B1(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__and3_1 _06629_ (.A(net857),
    .B(net848),
    .C(_00695_),
    .X(_00697_));
 sky130_fd_sc_hd__nor2_1 _06630_ (.A(_00696_),
    .B(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _06631_ (.A(net1550),
    .B(net860),
    .Y(_00699_));
 sky130_fd_sc_hd__and3_1 _06632_ (.A(net1496),
    .B(net1841),
    .C(_00699_),
    .X(_00700_));
 sky130_fd_sc_hd__xnor2_1 _06633_ (.A(_00698_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__a22oi_1 _06634_ (.A1(net1550),
    .A2(net1841),
    .B1(net860),
    .B2(net1496),
    .Y(_00702_));
 sky130_fd_sc_hd__and4_1 _06635_ (.A(net1496),
    .B(net1550),
    .C(net1841),
    .D(net860),
    .X(_00703_));
 sky130_fd_sc_hd__nor2_1 _06636_ (.A(_00702_),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__and3_1 _06637_ (.A(net1550),
    .B(net860),
    .C(net983),
    .X(_00705_));
 sky130_fd_sc_hd__a22o_1 _06638_ (.A1(net1550),
    .A2(net860),
    .B1(net983),
    .B2(net1496),
    .X(_00706_));
 sky130_fd_sc_hd__a21bo_1 _06639_ (.A1(net1496),
    .A2(_00705_),
    .B1_N(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__nand2_1 _06640_ (.A(net857),
    .B(net1841),
    .Y(_00708_));
 sky130_fd_sc_hd__a32o_1 _06641_ (.A1(net857),
    .A2(net1841),
    .A3(_00706_),
    .B1(_00705_),
    .B2(net1496),
    .X(_00709_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(_00704_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__or2_1 _06643_ (.A(_00704_),
    .B(_00709_),
    .X(_00711_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(_00710_),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__a22oi_1 _06645_ (.A1(net938),
    .A2(net848),
    .B1(net770),
    .B2(net857),
    .Y(_00713_));
 sky130_fd_sc_hd__or2_1 _06646_ (.A(_00694_),
    .B(_00713_),
    .X(_00714_));
 sky130_fd_sc_hd__or2_1 _06647_ (.A(_00712_),
    .B(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__a21o_1 _06648_ (.A1(_00710_),
    .A2(_00715_),
    .B1(_00701_),
    .X(_00716_));
 sky130_fd_sc_hd__nand3_1 _06649_ (.A(_00701_),
    .B(_00710_),
    .C(_00715_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(_00716_),
    .B(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand3_1 _06651_ (.A(_00694_),
    .B(_00716_),
    .C(_00717_),
    .Y(_00719_));
 sky130_fd_sc_hd__xor2_1 _06652_ (.A(_00694_),
    .B(_00718_),
    .X(_00720_));
 sky130_fd_sc_hd__xnor2_1 _06653_ (.A(_00712_),
    .B(_00714_),
    .Y(_00721_));
 sky130_fd_sc_hd__xnor2_1 _06654_ (.A(_00707_),
    .B(_00708_),
    .Y(_00722_));
 sky130_fd_sc_hd__and4_1 _06655_ (.A(net1550),
    .B(net857),
    .C(net860),
    .D(net983),
    .X(_00723_));
 sky130_fd_sc_hd__a22o_1 _06656_ (.A1(net857),
    .A2(net860),
    .B1(net983),
    .B2(net1550),
    .X(_00724_));
 sky130_fd_sc_hd__inv_2 _06657_ (.A(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__and4b_1 _06658_ (.A_N(_00723_),
    .B(_00724_),
    .C(net938),
    .D(net1841),
    .X(_00726_));
 sky130_fd_sc_hd__nor2_1 _06659_ (.A(_00723_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__or2_1 _06660_ (.A(_00722_),
    .B(_00727_),
    .X(_00728_));
 sky130_fd_sc_hd__xnor2_1 _06661_ (.A(_00722_),
    .B(_00727_),
    .Y(_00729_));
 sky130_fd_sc_hd__a22o_1 _06662_ (.A1(net878),
    .A2(net848),
    .B1(net770),
    .B2(net938),
    .X(_00730_));
 sky130_fd_sc_hd__inv_2 _06663_ (.A(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__and4_1 _06664_ (.A(net938),
    .B(net878),
    .C(net848),
    .D(net770),
    .X(_00732_));
 sky130_fd_sc_hd__or3_1 _06665_ (.A(_00729_),
    .B(_00731_),
    .C(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__a21o_1 _06666_ (.A1(_00728_),
    .A2(_00733_),
    .B1(_00721_),
    .X(_00734_));
 sky130_fd_sc_hd__nand3_1 _06667_ (.A(_00721_),
    .B(_00728_),
    .C(_00733_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand2_1 _06668_ (.A(_00734_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__inv_2 _06669_ (.A(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__nand2_1 _06670_ (.A(_00732_),
    .B(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__a21o_1 _06671_ (.A1(_00734_),
    .A2(_00738_),
    .B1(_00720_),
    .X(_00739_));
 sky130_fd_sc_hd__nand3_1 _06672_ (.A(_00720_),
    .B(_00734_),
    .C(_00738_),
    .Y(_00740_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(_00739_),
    .B(_00740_),
    .Y(_00741_));
 sky130_fd_sc_hd__xor2_1 _06674_ (.A(_00732_),
    .B(_00736_),
    .X(_00742_));
 sky130_fd_sc_hd__o21ai_1 _06675_ (.A1(_00731_),
    .A2(_00732_),
    .B1(_00729_),
    .Y(_00743_));
 sky130_fd_sc_hd__and2_1 _06676_ (.A(_00733_),
    .B(_00743_),
    .X(_00744_));
 sky130_fd_sc_hd__o2bb2a_1 _06677_ (.A1_N(net938),
    .A2_N(net1841),
    .B1(_00723_),
    .B2(_00725_),
    .X(_00745_));
 sky130_fd_sc_hd__or2_1 _06678_ (.A(_00726_),
    .B(_00745_),
    .X(_00746_));
 sky130_fd_sc_hd__and4_1 _06679_ (.A(net857),
    .B(net938),
    .C(net2522),
    .D(net983),
    .X(_00747_));
 sky130_fd_sc_hd__a22o_1 _06680_ (.A1(net938),
    .A2(net2522),
    .B1(net983),
    .B2(net857),
    .X(_00748_));
 sky130_fd_sc_hd__nand2b_1 _06681_ (.A_N(_00747_),
    .B(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _06682_ (.A(net878),
    .B(net1841),
    .Y(_00750_));
 sky130_fd_sc_hd__a31o_1 _06683_ (.A1(net878),
    .A2(net1841),
    .A3(_00748_),
    .B1(_00747_),
    .X(_00751_));
 sky130_fd_sc_hd__and2b_1 _06684_ (.A_N(_00746_),
    .B(_00751_),
    .X(_00752_));
 sky130_fd_sc_hd__xor2_1 _06685_ (.A(_00746_),
    .B(_00751_),
    .X(_00753_));
 sky130_fd_sc_hd__a22o_1 _06686_ (.A1(net803),
    .A2(net848),
    .B1(net770),
    .B2(net878),
    .X(_00754_));
 sky130_fd_sc_hd__and4_1 _06687_ (.A(net878),
    .B(net803),
    .C(net848),
    .D(net3720),
    .X(_00755_));
 sky130_fd_sc_hd__nand4_1 _06688_ (.A(net878),
    .B(net803),
    .C(net848),
    .D(net770),
    .Y(_00756_));
 sky130_fd_sc_hd__a22oi_1 _06689_ (.A1(net1496),
    .A2(net1729),
    .B1(_00754_),
    .B2(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hd__and4_1 _06690_ (.A(net1496),
    .B(net1729),
    .C(_00754_),
    .D(_00756_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _06691_ (.A(_00757_),
    .B(_00758_),
    .X(_00759_));
 sky130_fd_sc_hd__nor2_1 _06692_ (.A(_00753_),
    .B(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__o21ai_4 _06693_ (.A1(_00752_),
    .A2(_00760_),
    .B1(_00744_),
    .Y(_00761_));
 sky130_fd_sc_hd__or3_2 _06694_ (.A(_00744_),
    .B(_00752_),
    .C(_00760_),
    .X(_00762_));
 sky130_fd_sc_hd__o211ai_4 _06695_ (.A1(_00755_),
    .A2(_00758_),
    .B1(_00761_),
    .C1(_00762_),
    .Y(_00763_));
 sky130_fd_sc_hd__a21o_1 _06696_ (.A1(_00761_),
    .A2(_00763_),
    .B1(_00742_),
    .X(_00764_));
 sky130_fd_sc_hd__nor2_1 _06697_ (.A(_00741_),
    .B(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__and2_1 _06698_ (.A(_00741_),
    .B(_00764_),
    .X(_00766_));
 sky130_fd_sc_hd__nor2_1 _06699_ (.A(_00765_),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand3_1 _06700_ (.A(_00742_),
    .B(_00761_),
    .C(_00763_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _06701_ (.A(_00764_),
    .B(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__a211o_1 _06702_ (.A1(_00761_),
    .A2(_00762_),
    .B1(_00755_),
    .C1(_00758_),
    .X(_00770_));
 sky130_fd_sc_hd__xor2_1 _06703_ (.A(_00753_),
    .B(_00759_),
    .X(_00771_));
 sky130_fd_sc_hd__xnor2_1 _06704_ (.A(_00749_),
    .B(_00750_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand4_1 _06705_ (.A(net938),
    .B(net878),
    .C(net860),
    .D(net983),
    .Y(_00773_));
 sky130_fd_sc_hd__a22o_1 _06706_ (.A1(net878),
    .A2(net860),
    .B1(net983),
    .B2(net938),
    .X(_00774_));
 sky130_fd_sc_hd__and4_1 _06707_ (.A(net803),
    .B(net1841),
    .C(_00773_),
    .D(_00774_),
    .X(_00775_));
 sky130_fd_sc_hd__a41o_1 _06708_ (.A1(net938),
    .A2(net878),
    .A3(net860),
    .A4(net983),
    .B1(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__and2b_1 _06709_ (.A_N(_00772_),
    .B(_00776_),
    .X(_00777_));
 sky130_fd_sc_hd__nand4_1 _06710_ (.A(net803),
    .B(net806),
    .C(net848),
    .D(net770),
    .Y(_00778_));
 sky130_fd_sc_hd__a22o_1 _06711_ (.A1(net806),
    .A2(net2505),
    .B1(net770),
    .B2(net803),
    .X(_00779_));
 sky130_fd_sc_hd__nand2_1 _06712_ (.A(_00778_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _06713_ (.A(net1550),
    .B(net1729),
    .Y(_00781_));
 sky130_fd_sc_hd__xnor2_1 _06714_ (.A(_00780_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__xor2_1 _06715_ (.A(_00772_),
    .B(_00776_),
    .X(_00783_));
 sky130_fd_sc_hd__o21ba_1 _06716_ (.A1(_00782_),
    .A2(_00783_),
    .B1_N(_00777_),
    .X(_00784_));
 sky130_fd_sc_hd__and2b_1 _06717_ (.A_N(_00784_),
    .B(_00771_),
    .X(_00785_));
 sky130_fd_sc_hd__o21ai_1 _06718_ (.A1(_00780_),
    .A2(_00781_),
    .B1(_00778_),
    .Y(_00786_));
 sky130_fd_sc_hd__xnor2_1 _06719_ (.A(_00771_),
    .B(_00784_),
    .Y(_00787_));
 sky130_fd_sc_hd__and2_1 _06720_ (.A(_00786_),
    .B(_00787_),
    .X(_00788_));
 sky130_fd_sc_hd__o211ai_4 _06721_ (.A1(_00785_),
    .A2(_00788_),
    .B1(_00763_),
    .C1(_00770_),
    .Y(_00789_));
 sky130_fd_sc_hd__a211o_1 _06722_ (.A1(_00763_),
    .A2(_00770_),
    .B1(_00785_),
    .C1(_00788_),
    .X(_00790_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(_00789_),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__xnor2_1 _06724_ (.A(_00786_),
    .B(_00787_),
    .Y(_00792_));
 sky130_fd_sc_hd__xor2_1 _06725_ (.A(_00782_),
    .B(_00783_),
    .X(_00793_));
 sky130_fd_sc_hd__a22oi_1 _06726_ (.A1(net803),
    .A2(net1841),
    .B1(_00773_),
    .B2(_00774_),
    .Y(_00794_));
 sky130_fd_sc_hd__nor2_1 _06727_ (.A(_00775_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand4_1 _06728_ (.A(net878),
    .B(net803),
    .C(net2522),
    .D(net983),
    .Y(_00796_));
 sky130_fd_sc_hd__a22o_1 _06729_ (.A1(net803),
    .A2(net860),
    .B1(net983),
    .B2(net878),
    .X(_00797_));
 sky130_fd_sc_hd__nand4_1 _06730_ (.A(net806),
    .B(net1841),
    .C(_00796_),
    .D(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__and2_1 _06731_ (.A(_00796_),
    .B(_00798_),
    .X(_00799_));
 sky130_fd_sc_hd__and2b_1 _06732_ (.A_N(_00799_),
    .B(_00795_),
    .X(_00800_));
 sky130_fd_sc_hd__and4_1 _06733_ (.A(net806),
    .B(net1644),
    .C(net848),
    .D(net770),
    .X(_00801_));
 sky130_fd_sc_hd__a22o_1 _06734_ (.A1(net1644),
    .A2(net848),
    .B1(net770),
    .B2(net806),
    .X(_00802_));
 sky130_fd_sc_hd__inv_2 _06735_ (.A(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__and4b_1 _06736_ (.A_N(_00801_),
    .B(_00802_),
    .C(net857),
    .D(net1729),
    .X(_00804_));
 sky130_fd_sc_hd__o2bb2a_1 _06737_ (.A1_N(net857),
    .A2_N(net1729),
    .B1(_00801_),
    .B2(_00803_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _06738_ (.A(_00804_),
    .B(_00805_),
    .X(_00806_));
 sky130_fd_sc_hd__xnor2_1 _06739_ (.A(_00795_),
    .B(_00799_),
    .Y(_00807_));
 sky130_fd_sc_hd__and2b_1 _06740_ (.A_N(_00806_),
    .B(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__o21a_1 _06741_ (.A1(_00800_),
    .A2(_00808_),
    .B1(_00793_),
    .X(_00809_));
 sky130_fd_sc_hd__o211a_1 _06742_ (.A1(_00801_),
    .A2(_00804_),
    .B1(net1496),
    .C1(net764),
    .X(_00810_));
 sky130_fd_sc_hd__a211oi_1 _06743_ (.A1(net1496),
    .A2(net764),
    .B1(_00801_),
    .C1(_00804_),
    .Y(_00811_));
 sky130_fd_sc_hd__or2_1 _06744_ (.A(_00810_),
    .B(_00811_),
    .X(_00812_));
 sky130_fd_sc_hd__nor3_1 _06745_ (.A(_00793_),
    .B(_00800_),
    .C(_00808_),
    .Y(_00813_));
 sky130_fd_sc_hd__or3_1 _06746_ (.A(_00809_),
    .B(_00812_),
    .C(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__and2b_1 _06747_ (.A_N(_00809_),
    .B(_00814_),
    .X(_00815_));
 sky130_fd_sc_hd__nor2_1 _06748_ (.A(_00792_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__xor2_1 _06749_ (.A(_00792_),
    .B(_00815_),
    .X(_00817_));
 sky130_fd_sc_hd__and2_1 _06750_ (.A(_00810_),
    .B(_00817_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _06751_ (.A(_00816_),
    .B(_00818_),
    .X(_00819_));
 sky130_fd_sc_hd__and3_1 _06752_ (.A(_00789_),
    .B(_00790_),
    .C(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__o21bai_1 _06753_ (.A1(_00816_),
    .A2(_00818_),
    .B1_N(_00791_),
    .Y(_00821_));
 sky130_fd_sc_hd__a21oi_1 _06754_ (.A1(_00789_),
    .A2(_00821_),
    .B1(_00769_),
    .Y(_00822_));
 sky130_fd_sc_hd__xor2_2 _06755_ (.A(_00769_),
    .B(_00789_),
    .X(_00823_));
 sky130_fd_sc_hd__xnor2_2 _06756_ (.A(_00791_),
    .B(_00819_),
    .Y(_00824_));
 sky130_fd_sc_hd__xnor2_1 _06757_ (.A(_00810_),
    .B(_00817_),
    .Y(_00825_));
 sky130_fd_sc_hd__o21ai_1 _06758_ (.A1(_00809_),
    .A2(_00813_),
    .B1(_00812_),
    .Y(_00826_));
 sky130_fd_sc_hd__xnor2_1 _06759_ (.A(_00806_),
    .B(_00807_),
    .Y(_00827_));
 sky130_fd_sc_hd__a22o_1 _06760_ (.A1(net806),
    .A2(net1841),
    .B1(_00796_),
    .B2(_00797_),
    .X(_00828_));
 sky130_fd_sc_hd__nand4_1 _06761_ (.A(net803),
    .B(net806),
    .C(net860),
    .D(net983),
    .Y(_00829_));
 sky130_fd_sc_hd__and2_1 _06762_ (.A(net1644),
    .B(net1841),
    .X(_00830_));
 sky130_fd_sc_hd__a22o_1 _06763_ (.A1(net806),
    .A2(net860),
    .B1(net983),
    .B2(net803),
    .X(_00831_));
 sky130_fd_sc_hd__nand3_1 _06764_ (.A(_00829_),
    .B(_00830_),
    .C(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__a21bo_1 _06765_ (.A1(_00830_),
    .A2(_00831_),
    .B1_N(_00829_),
    .X(_00833_));
 sky130_fd_sc_hd__nand3_1 _06766_ (.A(_00798_),
    .B(_00828_),
    .C(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__and4_1 _06767_ (.A(net938),
    .B(net1644),
    .C(net770),
    .D(net1729),
    .X(_00835_));
 sky130_fd_sc_hd__a22oi_1 _06768_ (.A1(net1644),
    .A2(net770),
    .B1(net1729),
    .B2(net938),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2_1 _06769_ (.A(_00835_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__a21o_1 _06770_ (.A1(_00798_),
    .A2(_00828_),
    .B1(_00833_),
    .X(_00838_));
 sky130_fd_sc_hd__nand3_1 _06771_ (.A(_00834_),
    .B(_00837_),
    .C(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__and2_1 _06772_ (.A(_00834_),
    .B(_00839_),
    .X(_00840_));
 sky130_fd_sc_hd__and2b_1 _06773_ (.A_N(_00840_),
    .B(_00827_),
    .X(_00841_));
 sky130_fd_sc_hd__a21o_1 _06774_ (.A1(net1550),
    .A2(net764),
    .B1(_00835_),
    .X(_00842_));
 sky130_fd_sc_hd__nand3_1 _06775_ (.A(net1550),
    .B(net764),
    .C(_00835_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(_00842_),
    .B(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(net1496),
    .B(net2041),
    .Y(_00845_));
 sky130_fd_sc_hd__xor2_1 _06778_ (.A(_00844_),
    .B(_00845_),
    .X(_00846_));
 sky130_fd_sc_hd__xnor2_1 _06779_ (.A(_00827_),
    .B(_00840_),
    .Y(_00847_));
 sky130_fd_sc_hd__and2_1 _06780_ (.A(_00846_),
    .B(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__o211a_1 _06781_ (.A1(_00841_),
    .A2(_00848_),
    .B1(_00814_),
    .C1(_00826_),
    .X(_00849_));
 sky130_fd_sc_hd__o21a_1 _06782_ (.A1(_00844_),
    .A2(_00845_),
    .B1(_00843_),
    .X(_00850_));
 sky130_fd_sc_hd__a211oi_1 _06783_ (.A1(_00814_),
    .A2(_00826_),
    .B1(_00841_),
    .C1(_00848_),
    .Y(_00851_));
 sky130_fd_sc_hd__nor2_1 _06784_ (.A(_00849_),
    .B(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hd__o21bai_1 _06785_ (.A1(_00850_),
    .A2(_00851_),
    .B1_N(_00849_),
    .Y(_00853_));
 sky130_fd_sc_hd__and2b_1 _06786_ (.A_N(_00853_),
    .B(_00825_),
    .X(_00854_));
 sky130_fd_sc_hd__nand2b_1 _06787_ (.A_N(_00853_),
    .B(_00825_),
    .Y(_00855_));
 sky130_fd_sc_hd__and2b_1 _06788_ (.A_N(_00825_),
    .B(_00853_),
    .X(_00856_));
 sky130_fd_sc_hd__xnor2_2 _06789_ (.A(_00850_),
    .B(_00852_),
    .Y(_00857_));
 sky130_fd_sc_hd__xor2_1 _06790_ (.A(_00846_),
    .B(_00847_),
    .X(_00858_));
 sky130_fd_sc_hd__a21o_1 _06791_ (.A1(_00834_),
    .A2(_00838_),
    .B1(_00837_),
    .X(_00859_));
 sky130_fd_sc_hd__a21o_1 _06792_ (.A1(_00829_),
    .A2(_00831_),
    .B1(_00830_),
    .X(_00860_));
 sky130_fd_sc_hd__and4_1 _06793_ (.A(net806),
    .B(net1644),
    .C(net860),
    .D(net983),
    .X(_00861_));
 sky130_fd_sc_hd__and3_1 _06794_ (.A(_00832_),
    .B(_00860_),
    .C(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(net878),
    .B(net1729),
    .Y(_00863_));
 sky130_fd_sc_hd__a21oi_1 _06796_ (.A1(_00832_),
    .A2(_00860_),
    .B1(_00861_),
    .Y(_00864_));
 sky130_fd_sc_hd__or3_1 _06797_ (.A(_00862_),
    .B(_00863_),
    .C(_00864_),
    .X(_00865_));
 sky130_fd_sc_hd__o21bai_1 _06798_ (.A1(_00863_),
    .A2(_00864_),
    .B1_N(_00862_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand3_2 _06799_ (.A(_00839_),
    .B(_00859_),
    .C(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__a22o_1 _06800_ (.A1(net857),
    .A2(net764),
    .B1(net2041),
    .B2(net1550),
    .X(_00868_));
 sky130_fd_sc_hd__nand4_2 _06801_ (.A(net1550),
    .B(net2584),
    .C(net764),
    .D(net2041),
    .Y(_00869_));
 sky130_fd_sc_hd__and2_1 _06802_ (.A(_00868_),
    .B(_00869_),
    .X(_00870_));
 sky130_fd_sc_hd__a21o_1 _06803_ (.A1(_00839_),
    .A2(_00859_),
    .B1(_00866_),
    .X(_00871_));
 sky130_fd_sc_hd__nand3_2 _06804_ (.A(_00867_),
    .B(_00870_),
    .C(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_1 _06805_ (.A(_00867_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _06806_ (.A(_00858_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__xnor2_1 _06807_ (.A(_00858_),
    .B(_00873_),
    .Y(_00875_));
 sky130_fd_sc_hd__o21ai_2 _06808_ (.A1(_00869_),
    .A2(_00875_),
    .B1(_00874_),
    .Y(_00876_));
 sky130_fd_sc_hd__and2_1 _06809_ (.A(_00857_),
    .B(_00876_),
    .X(_00877_));
 sky130_fd_sc_hd__xnor2_1 _06810_ (.A(_00869_),
    .B(_00875_),
    .Y(_00878_));
 sky130_fd_sc_hd__a21o_1 _06811_ (.A1(_00867_),
    .A2(_00871_),
    .B1(_00870_),
    .X(_00879_));
 sky130_fd_sc_hd__o21ai_1 _06812_ (.A1(_00862_),
    .A2(_00864_),
    .B1(_00863_),
    .Y(_00880_));
 sky130_fd_sc_hd__a22oi_1 _06813_ (.A1(net1644),
    .A2(net860),
    .B1(net983),
    .B2(net806),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2_1 _06814_ (.A(_00861_),
    .B(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _06815_ (.A(net803),
    .B(net1729),
    .Y(_00883_));
 sky130_fd_sc_hd__and3_1 _06816_ (.A(net803),
    .B(net1729),
    .C(_00882_),
    .X(_00884_));
 sky130_fd_sc_hd__nand3_1 _06817_ (.A(_00865_),
    .B(_00880_),
    .C(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__a22oi_1 _06818_ (.A1(net938),
    .A2(net764),
    .B1(net2041),
    .B2(net857),
    .Y(_00886_));
 sky130_fd_sc_hd__and4_1 _06819_ (.A(net2582),
    .B(net938),
    .C(net3725),
    .D(net2041),
    .X(_00887_));
 sky130_fd_sc_hd__nor2_1 _06820_ (.A(_00886_),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a21o_1 _06821_ (.A1(_00865_),
    .A2(_00880_),
    .B1(_00884_),
    .X(_00889_));
 sky130_fd_sc_hd__nand3_1 _06822_ (.A(_00885_),
    .B(_00888_),
    .C(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__a21bo_1 _06823_ (.A1(_00888_),
    .A2(_00889_),
    .B1_N(_00885_),
    .X(_00891_));
 sky130_fd_sc_hd__nand3_2 _06824_ (.A(_00872_),
    .B(_00879_),
    .C(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__a21o_1 _06825_ (.A1(_00872_),
    .A2(_00879_),
    .B1(_00891_),
    .X(_00893_));
 sky130_fd_sc_hd__nand3_2 _06826_ (.A(_00887_),
    .B(_00892_),
    .C(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__a21o_1 _06827_ (.A1(_00892_),
    .A2(_00894_),
    .B1(_00878_),
    .X(_00895_));
 sky130_fd_sc_hd__inv_2 _06828_ (.A(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__and3_1 _06829_ (.A(_00878_),
    .B(_00892_),
    .C(_00894_),
    .X(_00897_));
 sky130_fd_sc_hd__a21o_1 _06830_ (.A1(_00892_),
    .A2(_00893_),
    .B1(_00887_),
    .X(_00898_));
 sky130_fd_sc_hd__a21o_1 _06831_ (.A1(_00885_),
    .A2(_00889_),
    .B1(_00888_),
    .X(_00899_));
 sky130_fd_sc_hd__xnor2_1 _06832_ (.A(_00882_),
    .B(_00883_),
    .Y(_00900_));
 sky130_fd_sc_hd__and4_1 _06833_ (.A(net806),
    .B(net1644),
    .C(net3643),
    .D(net1729),
    .X(_00901_));
 sky130_fd_sc_hd__inv_2 _06834_ (.A(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_00900_),
    .B(_00901_),
    .Y(_00903_));
 sky130_fd_sc_hd__a22oi_1 _06836_ (.A1(net878),
    .A2(net764),
    .B1(net2041),
    .B2(net3646),
    .Y(_00904_));
 sky130_fd_sc_hd__and4_1 _06837_ (.A(net3646),
    .B(net878),
    .C(net764),
    .D(net2041),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _06838_ (.A(_00904_),
    .B(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_2 _06839_ (.A(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__xnor2_1 _06840_ (.A(_00900_),
    .B(_00901_),
    .Y(_00908_));
 sky130_fd_sc_hd__o21ai_1 _06841_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00903_),
    .Y(_00909_));
 sky130_fd_sc_hd__and3_1 _06842_ (.A(_00890_),
    .B(_00899_),
    .C(_00909_),
    .X(_00910_));
 sky130_fd_sc_hd__a21o_1 _06843_ (.A1(_00890_),
    .A2(_00899_),
    .B1(_00909_),
    .X(_00911_));
 sky130_fd_sc_hd__and2b_1 _06844_ (.A_N(_00910_),
    .B(_00911_),
    .X(_00912_));
 sky130_fd_sc_hd__a21o_1 _06845_ (.A1(_00905_),
    .A2(_00911_),
    .B1(_00910_),
    .X(_00913_));
 sky130_fd_sc_hd__and3_1 _06846_ (.A(_00894_),
    .B(_00898_),
    .C(_00913_),
    .X(_00914_));
 sky130_fd_sc_hd__nand3_1 _06847_ (.A(_00894_),
    .B(_00898_),
    .C(_00913_),
    .Y(_00915_));
 sky130_fd_sc_hd__a21oi_1 _06848_ (.A1(_00894_),
    .A2(_00898_),
    .B1(_00913_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _06849_ (.A(_00914_),
    .B(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__xnor2_1 _06850_ (.A(_00905_),
    .B(_00912_),
    .Y(_00918_));
 sky130_fd_sc_hd__xnor2_1 _06851_ (.A(_00906_),
    .B(_00908_),
    .Y(_00919_));
 sky130_fd_sc_hd__and4_1 _06852_ (.A(net3651),
    .B(net803),
    .C(net764),
    .D(net2041),
    .X(_00920_));
 sky130_fd_sc_hd__inv_2 _06853_ (.A(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__a22o_1 _06854_ (.A1(net1644),
    .A2(net3643),
    .B1(net1729),
    .B2(net806),
    .X(_00922_));
 sky130_fd_sc_hd__a22o_1 _06855_ (.A1(net803),
    .A2(net764),
    .B1(net2041),
    .B2(net3651),
    .X(_00923_));
 sky130_fd_sc_hd__or4bb_2 _06856_ (.A(_00901_),
    .B(_00920_),
    .C_N(_00922_),
    .D_N(_00923_),
    .X(_00924_));
 sky130_fd_sc_hd__a21boi_1 _06857_ (.A1(_00921_),
    .A2(_00924_),
    .B1_N(_00919_),
    .Y(_00925_));
 sky130_fd_sc_hd__and3b_1 _06858_ (.A_N(_00919_),
    .B(_00921_),
    .C(_00924_),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_1 _06859_ (.A1(_00902_),
    .A2(_00922_),
    .B1(_00923_),
    .B2(_00921_),
    .X(_00927_));
 sky130_fd_sc_hd__and4_2 _06860_ (.A(net2203),
    .B(net806),
    .C(net764),
    .D(net2041),
    .X(_00928_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(net1644),
    .B(net1729),
    .Y(_00929_));
 sky130_fd_sc_hd__a22o_1 _06862_ (.A1(net2054),
    .A2(net764),
    .B1(net2041),
    .B2(net2203),
    .X(_00930_));
 sky130_fd_sc_hd__inv_2 _06863_ (.A(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__nor3_1 _06864_ (.A(_00928_),
    .B(_00929_),
    .C(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__or3_1 _06865_ (.A(_00928_),
    .B(_00929_),
    .C(_00931_),
    .X(_00933_));
 sky130_fd_sc_hd__o211ai_2 _06866_ (.A1(_00928_),
    .A2(_00932_),
    .B1(_00924_),
    .C1(_00927_),
    .Y(_00934_));
 sky130_fd_sc_hd__o21ai_1 _06867_ (.A1(_00928_),
    .A2(_00931_),
    .B1(_00929_),
    .Y(_00935_));
 sky130_fd_sc_hd__and4_1 _06868_ (.A(net806),
    .B(net1644),
    .C(net764),
    .D(net2041),
    .X(_00936_));
 sky130_fd_sc_hd__and3_1 _06869_ (.A(_00933_),
    .B(_00935_),
    .C(_00936_),
    .X(_00937_));
 sky130_fd_sc_hd__a211o_1 _06870_ (.A1(_00924_),
    .A2(_00927_),
    .B1(_00928_),
    .C1(_00932_),
    .X(_00938_));
 sky130_fd_sc_hd__and2_1 _06871_ (.A(_00934_),
    .B(_00938_),
    .X(_00939_));
 sky130_fd_sc_hd__nand2_1 _06872_ (.A(_00937_),
    .B(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__a211oi_2 _06873_ (.A1(_00934_),
    .A2(_00940_),
    .B1(_00925_),
    .C1(_00926_),
    .Y(_00941_));
 sky130_fd_sc_hd__or2_1 _06874_ (.A(_00925_),
    .B(_00941_),
    .X(_00942_));
 sky130_fd_sc_hd__inv_2 _06875_ (.A(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__nor2_1 _06876_ (.A(_00918_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__o31a_1 _06877_ (.A1(_00916_),
    .A2(_00918_),
    .A3(_00943_),
    .B1(_00915_),
    .X(_00945_));
 sky130_fd_sc_hd__o21ai_4 _06878_ (.A1(_00897_),
    .A2(_00945_),
    .B1(_00895_),
    .Y(_00946_));
 sky130_fd_sc_hd__xor2_2 _06879_ (.A(_00857_),
    .B(_00876_),
    .X(_00947_));
 sky130_fd_sc_hd__a21o_1 _06880_ (.A1(_00946_),
    .A2(_00947_),
    .B1(_00877_),
    .X(_00948_));
 sky130_fd_sc_hd__a211o_1 _06881_ (.A1(_00946_),
    .A2(_00947_),
    .B1(_00856_),
    .C1(_00877_),
    .X(_00949_));
 sky130_fd_sc_hd__nand2_1 _06882_ (.A(_00855_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__a41o_1 _06883_ (.A1(_00823_),
    .A2(_00824_),
    .A3(_00855_),
    .A4(_00949_),
    .B1(_00822_),
    .X(_00951_));
 sky130_fd_sc_hd__xor2_1 _06884_ (.A(_00767_),
    .B(_00951_),
    .X(_00952_));
 sky130_fd_sc_hd__a22oi_1 _06885_ (.A1(net697),
    .A2(net2152),
    .B1(net995),
    .B2(net1456),
    .Y(_00953_));
 sky130_fd_sc_hd__and4_1 _06886_ (.A(net1456),
    .B(net697),
    .C(net2152),
    .D(net995),
    .X(_00954_));
 sky130_fd_sc_hd__or2_1 _06887_ (.A(_00953_),
    .B(_00954_),
    .X(_00955_));
 sky130_fd_sc_hd__nand2_1 _06888_ (.A(net697),
    .B(net995),
    .Y(_00956_));
 sky130_fd_sc_hd__and4_1 _06889_ (.A(net1456),
    .B(net697),
    .C(net995),
    .D(net842),
    .X(_00957_));
 sky130_fd_sc_hd__a22o_1 _06890_ (.A1(net697),
    .A2(net995),
    .B1(net842),
    .B2(net1456),
    .X(_00958_));
 sky130_fd_sc_hd__and2b_1 _06891_ (.A_N(_00957_),
    .B(_00958_),
    .X(_00959_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(net776),
    .B(net2152),
    .Y(_00960_));
 sky130_fd_sc_hd__a31oi_2 _06893_ (.A1(net776),
    .A2(net2152),
    .A3(_00958_),
    .B1(_00957_),
    .Y(_00961_));
 sky130_fd_sc_hd__xor2_1 _06894_ (.A(_00955_),
    .B(_00961_),
    .X(_00962_));
 sky130_fd_sc_hd__and3_1 _06895_ (.A(net776),
    .B(net752),
    .C(_00962_),
    .X(_00963_));
 sky130_fd_sc_hd__a21oi_1 _06896_ (.A1(net776),
    .A2(net752),
    .B1(_00962_),
    .Y(_00964_));
 sky130_fd_sc_hd__or2_1 _06897_ (.A(_00963_),
    .B(_00964_),
    .X(_00965_));
 sky130_fd_sc_hd__xnor2_1 _06898_ (.A(_00959_),
    .B(_00960_),
    .Y(_00966_));
 sky130_fd_sc_hd__and4_1 _06899_ (.A(net697),
    .B(net776),
    .C(net995),
    .D(net842),
    .X(_00967_));
 sky130_fd_sc_hd__a22o_1 _06900_ (.A1(net776),
    .A2(net995),
    .B1(net842),
    .B2(net697),
    .X(_00968_));
 sky130_fd_sc_hd__inv_2 _06901_ (.A(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__and4b_1 _06902_ (.A_N(_00967_),
    .B(_00968_),
    .C(net833),
    .D(net2152),
    .X(_00970_));
 sky130_fd_sc_hd__or2_1 _06903_ (.A(_00967_),
    .B(_00970_),
    .X(_00971_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_00966_),
    .B(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__xor2_1 _06905_ (.A(_00966_),
    .B(_00971_),
    .X(_00973_));
 sky130_fd_sc_hd__nand3_1 _06906_ (.A(net833),
    .B(net752),
    .C(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__a21oi_1 _06907_ (.A1(_00972_),
    .A2(_00974_),
    .B1(_00965_),
    .Y(_00975_));
 sky130_fd_sc_hd__and3_1 _06908_ (.A(_00965_),
    .B(_00972_),
    .C(_00974_),
    .X(_00976_));
 sky130_fd_sc_hd__nor2_1 _06909_ (.A(_00975_),
    .B(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__a21o_1 _06910_ (.A1(net833),
    .A2(net752),
    .B1(_00973_),
    .X(_00978_));
 sky130_fd_sc_hd__and2_1 _06911_ (.A(_00974_),
    .B(_00978_),
    .X(_00979_));
 sky130_fd_sc_hd__o2bb2a_1 _06912_ (.A1_N(net833),
    .A2_N(net2152),
    .B1(_00967_),
    .B2(_00969_),
    .X(_00980_));
 sky130_fd_sc_hd__or2_1 _06913_ (.A(_00970_),
    .B(_00980_),
    .X(_00981_));
 sky130_fd_sc_hd__and4_1 _06914_ (.A(net776),
    .B(net833),
    .C(net995),
    .D(net842),
    .X(_00982_));
 sky130_fd_sc_hd__a22o_1 _06915_ (.A1(net833),
    .A2(net995),
    .B1(net842),
    .B2(net776),
    .X(_00983_));
 sky130_fd_sc_hd__nand2b_1 _06916_ (.A_N(_00982_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _06917_ (.A(net800),
    .B(net2152),
    .Y(_00985_));
 sky130_fd_sc_hd__a31o_1 _06918_ (.A1(net800),
    .A2(net2152),
    .A3(_00983_),
    .B1(_00982_),
    .X(_00986_));
 sky130_fd_sc_hd__and2b_1 _06919_ (.A_N(_00981_),
    .B(_00986_),
    .X(_00987_));
 sky130_fd_sc_hd__xor2_2 _06920_ (.A(_00981_),
    .B(_00986_),
    .X(_00988_));
 sky130_fd_sc_hd__a22oi_1 _06921_ (.A1(net800),
    .A2(net752),
    .B1(net926),
    .B2(net1456),
    .Y(_00989_));
 sky130_fd_sc_hd__and4_2 _06922_ (.A(net1456),
    .B(net800),
    .C(net752),
    .D(net926),
    .X(_00990_));
 sky130_fd_sc_hd__nor2_1 _06923_ (.A(_00989_),
    .B(_00990_),
    .Y(_00991_));
 sky130_fd_sc_hd__and2b_1 _06924_ (.A_N(_00988_),
    .B(_00991_),
    .X(_00992_));
 sky130_fd_sc_hd__o21a_1 _06925_ (.A1(_00987_),
    .A2(_00992_),
    .B1(_00979_),
    .X(_00993_));
 sky130_fd_sc_hd__nor3_1 _06926_ (.A(_00979_),
    .B(_00987_),
    .C(_00992_),
    .Y(_00994_));
 sky130_fd_sc_hd__nor2_2 _06927_ (.A(_00993_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__a21o_1 _06928_ (.A1(_00990_),
    .A2(_00995_),
    .B1(_00993_),
    .X(_00996_));
 sky130_fd_sc_hd__and2_1 _06929_ (.A(_00977_),
    .B(_00996_),
    .X(_00997_));
 sky130_fd_sc_hd__xnor2_1 _06930_ (.A(_00977_),
    .B(_00996_),
    .Y(_00998_));
 sky130_fd_sc_hd__xnor2_4 _06931_ (.A(_00990_),
    .B(_00995_),
    .Y(_00999_));
 sky130_fd_sc_hd__xnor2_2 _06932_ (.A(_00988_),
    .B(_00991_),
    .Y(_01000_));
 sky130_fd_sc_hd__xnor2_1 _06933_ (.A(_00984_),
    .B(_00985_),
    .Y(_01001_));
 sky130_fd_sc_hd__and4_1 _06934_ (.A(net833),
    .B(net800),
    .C(net995),
    .D(net842),
    .X(_01002_));
 sky130_fd_sc_hd__a22o_1 _06935_ (.A1(net800),
    .A2(net995),
    .B1(net842),
    .B2(net833),
    .X(_01003_));
 sky130_fd_sc_hd__nand2b_1 _06936_ (.A_N(_01002_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand2_1 _06937_ (.A(net929),
    .B(net2152),
    .Y(_01005_));
 sky130_fd_sc_hd__a31o_1 _06938_ (.A1(net929),
    .A2(net2152),
    .A3(_01003_),
    .B1(_01002_),
    .X(_01006_));
 sky130_fd_sc_hd__and2b_1 _06939_ (.A_N(_01001_),
    .B(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__xor2_1 _06940_ (.A(_01001_),
    .B(_01006_),
    .X(_01008_));
 sky130_fd_sc_hd__a22o_1 _06941_ (.A1(net929),
    .A2(net752),
    .B1(net926),
    .B2(net697),
    .X(_01009_));
 sky130_fd_sc_hd__and4_1 _06942_ (.A(net697),
    .B(net929),
    .C(net752),
    .D(net926),
    .X(_01010_));
 sky130_fd_sc_hd__nand4_1 _06943_ (.A(net697),
    .B(net929),
    .C(net752),
    .D(net926),
    .Y(_01011_));
 sky130_fd_sc_hd__a22oi_1 _06944_ (.A1(net1456),
    .A2(net998),
    .B1(_01009_),
    .B2(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__and4_1 _06945_ (.A(net1456),
    .B(net998),
    .C(_01009_),
    .D(_01011_),
    .X(_01013_));
 sky130_fd_sc_hd__or2_1 _06946_ (.A(_01012_),
    .B(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2_1 _06947_ (.A(_01008_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__o21ai_4 _06948_ (.A1(_01007_),
    .A2(_01015_),
    .B1(_01000_),
    .Y(_01016_));
 sky130_fd_sc_hd__or3_2 _06949_ (.A(_01000_),
    .B(_01007_),
    .C(_01015_),
    .X(_01017_));
 sky130_fd_sc_hd__o211ai_4 _06950_ (.A1(_01010_),
    .A2(_01013_),
    .B1(_01016_),
    .C1(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_2 _06951_ (.A(_01016_),
    .B(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2b_1 _06952_ (.A_N(_00999_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__nor2_1 _06953_ (.A(_00998_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(_00998_),
    .B(_01020_),
    .Y(_01022_));
 sky130_fd_sc_hd__and2b_1 _06955_ (.A_N(_01021_),
    .B(_01022_),
    .X(_01023_));
 sky130_fd_sc_hd__xor2_4 _06956_ (.A(_00999_),
    .B(_01019_),
    .X(_01024_));
 sky130_fd_sc_hd__a211o_1 _06957_ (.A1(_01016_),
    .A2(_01017_),
    .B1(_01010_),
    .C1(_01013_),
    .X(_01025_));
 sky130_fd_sc_hd__xor2_1 _06958_ (.A(_01008_),
    .B(_01014_),
    .X(_01026_));
 sky130_fd_sc_hd__xnor2_2 _06959_ (.A(_01004_),
    .B(_01005_),
    .Y(_01027_));
 sky130_fd_sc_hd__nand4_2 _06960_ (.A(net800),
    .B(net929),
    .C(net995),
    .D(net842),
    .Y(_01028_));
 sky130_fd_sc_hd__a22o_1 _06961_ (.A1(net929),
    .A2(net995),
    .B1(net842),
    .B2(net800),
    .X(_01029_));
 sky130_fd_sc_hd__nand4_2 _06962_ (.A(net911),
    .B(net2152),
    .C(_01028_),
    .D(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_1 _06963_ (.A(_01028_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__and2b_1 _06964_ (.A_N(_01027_),
    .B(_01031_),
    .X(_01032_));
 sky130_fd_sc_hd__nand4_2 _06965_ (.A(net776),
    .B(net911),
    .C(net752),
    .D(net926),
    .Y(_01033_));
 sky130_fd_sc_hd__a22o_1 _06966_ (.A1(net911),
    .A2(net2768),
    .B1(net926),
    .B2(net776),
    .X(_01034_));
 sky130_fd_sc_hd__nand2_2 _06967_ (.A(_01033_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_1 _06968_ (.A(net697),
    .B(net998),
    .Y(_01036_));
 sky130_fd_sc_hd__xnor2_2 _06969_ (.A(_01035_),
    .B(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__xor2_2 _06970_ (.A(_01027_),
    .B(_01031_),
    .X(_01038_));
 sky130_fd_sc_hd__nor2_1 _06971_ (.A(_01037_),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__o21a_1 _06972_ (.A1(_01032_),
    .A2(_01039_),
    .B1(_01026_),
    .X(_01040_));
 sky130_fd_sc_hd__o21ai_2 _06973_ (.A1(_01035_),
    .A2(_01036_),
    .B1(_01033_),
    .Y(_01041_));
 sky130_fd_sc_hd__or3_1 _06974_ (.A(_01026_),
    .B(_01032_),
    .C(_01039_),
    .X(_01042_));
 sky130_fd_sc_hd__nand2b_1 _06975_ (.A_N(_01040_),
    .B(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__and2b_1 _06976_ (.A_N(_01043_),
    .B(_01041_),
    .X(_01044_));
 sky130_fd_sc_hd__o211ai_2 _06977_ (.A1(_01040_),
    .A2(_01044_),
    .B1(_01018_),
    .C1(_01025_),
    .Y(_01045_));
 sky130_fd_sc_hd__inv_2 _06978_ (.A(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__a211o_1 _06979_ (.A1(_01018_),
    .A2(_01025_),
    .B1(_01040_),
    .C1(_01044_),
    .X(_01047_));
 sky130_fd_sc_hd__nand2_2 _06980_ (.A(_01045_),
    .B(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__xnor2_2 _06981_ (.A(_01041_),
    .B(_01043_),
    .Y(_01049_));
 sky130_fd_sc_hd__xor2_2 _06982_ (.A(_01037_),
    .B(_01038_),
    .X(_01050_));
 sky130_fd_sc_hd__a22o_1 _06983_ (.A1(net911),
    .A2(net2152),
    .B1(_01028_),
    .B2(_01029_),
    .X(_01051_));
 sky130_fd_sc_hd__nand4_1 _06984_ (.A(net929),
    .B(net911),
    .C(net995),
    .D(net842),
    .Y(_01052_));
 sky130_fd_sc_hd__and2_1 _06985_ (.A(net88),
    .B(net2152),
    .X(_01053_));
 sky130_fd_sc_hd__a22o_1 _06986_ (.A1(net911),
    .A2(net995),
    .B1(net2343),
    .B2(net929),
    .X(_01054_));
 sky130_fd_sc_hd__nand3_1 _06987_ (.A(_01052_),
    .B(_01053_),
    .C(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__a21bo_1 _06988_ (.A1(_01053_),
    .A2(_01054_),
    .B1_N(_01052_),
    .X(_01056_));
 sky130_fd_sc_hd__nand3_1 _06989_ (.A(_01030_),
    .B(_01051_),
    .C(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__and4_1 _06990_ (.A(net833),
    .B(net88),
    .C(net752),
    .D(net926),
    .X(_01058_));
 sky130_fd_sc_hd__a22o_1 _06991_ (.A1(net88),
    .A2(net752),
    .B1(net926),
    .B2(net833),
    .X(_01059_));
 sky130_fd_sc_hd__and2b_1 _06992_ (.A_N(_01058_),
    .B(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(net776),
    .B(net998),
    .Y(_01061_));
 sky130_fd_sc_hd__xnor2_1 _06994_ (.A(_01060_),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__a21o_1 _06995_ (.A1(_01030_),
    .A2(_01051_),
    .B1(_01056_),
    .X(_01063_));
 sky130_fd_sc_hd__nand3_1 _06996_ (.A(_01057_),
    .B(_01062_),
    .C(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__and2_1 _06997_ (.A(_01057_),
    .B(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__and2b_1 _06998_ (.A_N(_01065_),
    .B(_01050_),
    .X(_01066_));
 sky130_fd_sc_hd__a31oi_2 _06999_ (.A1(net776),
    .A2(net998),
    .A3(_01059_),
    .B1(_01058_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(net1456),
    .B(net153),
    .Y(_01068_));
 sky130_fd_sc_hd__nor2_1 _07001_ (.A(_01067_),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__xnor2_1 _07002_ (.A(_01067_),
    .B(_01068_),
    .Y(_01070_));
 sky130_fd_sc_hd__and2b_1 _07003_ (.A_N(_01050_),
    .B(_01065_),
    .X(_01071_));
 sky130_fd_sc_hd__xnor2_1 _07004_ (.A(_01050_),
    .B(_01065_),
    .Y(_01072_));
 sky130_fd_sc_hd__o21bai_2 _07005_ (.A1(_01070_),
    .A2(_01071_),
    .B1_N(_01066_),
    .Y(_01073_));
 sky130_fd_sc_hd__and2_1 _07006_ (.A(_01049_),
    .B(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__xor2_2 _07007_ (.A(_01049_),
    .B(_01073_),
    .X(_01075_));
 sky130_fd_sc_hd__and2_1 _07008_ (.A(_01069_),
    .B(_01075_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_2 _07009_ (.A(_01074_),
    .B(_01076_),
    .X(_01077_));
 sky130_fd_sc_hd__o21ba_1 _07010_ (.A1(_01074_),
    .A2(_01076_),
    .B1_N(_01048_),
    .X(_01078_));
 sky130_fd_sc_hd__o21ba_1 _07011_ (.A1(_01046_),
    .A2(_01078_),
    .B1_N(_01024_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_4 _07012_ (.A(_01024_),
    .B(_01046_),
    .Y(_01080_));
 sky130_fd_sc_hd__xnor2_4 _07013_ (.A(_01048_),
    .B(_01077_),
    .Y(_01081_));
 sky130_fd_sc_hd__xnor2_2 _07014_ (.A(_01069_),
    .B(_01075_),
    .Y(_01082_));
 sky130_fd_sc_hd__xnor2_1 _07015_ (.A(_01070_),
    .B(_01072_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21o_1 _07016_ (.A1(_01057_),
    .A2(_01063_),
    .B1(_01062_),
    .X(_01084_));
 sky130_fd_sc_hd__a21o_1 _07017_ (.A1(_01052_),
    .A2(_01054_),
    .B1(_01053_),
    .X(_01085_));
 sky130_fd_sc_hd__and4_1 _07018_ (.A(net911),
    .B(net88),
    .C(net2349),
    .D(net2343),
    .X(_01086_));
 sky130_fd_sc_hd__nand4_1 _07019_ (.A(net911),
    .B(net88),
    .C(net2349),
    .D(net842),
    .Y(_01087_));
 sky130_fd_sc_hd__nand3_1 _07020_ (.A(_01055_),
    .B(_01085_),
    .C(_01086_),
    .Y(_01088_));
 sky130_fd_sc_hd__a22oi_1 _07021_ (.A1(net800),
    .A2(net926),
    .B1(net998),
    .B2(net833),
    .Y(_01089_));
 sky130_fd_sc_hd__and4_1 _07022_ (.A(net833),
    .B(net800),
    .C(net926),
    .D(net2068),
    .X(_01090_));
 sky130_fd_sc_hd__nor2_1 _07023_ (.A(_01089_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__a21o_1 _07024_ (.A1(_01055_),
    .A2(_01085_),
    .B1(_01086_),
    .X(_01092_));
 sky130_fd_sc_hd__nand3_1 _07025_ (.A(_01088_),
    .B(_01091_),
    .C(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__a21bo_1 _07026_ (.A1(_01091_),
    .A2(_01092_),
    .B1_N(_01088_),
    .X(_01094_));
 sky130_fd_sc_hd__nand3_1 _07027_ (.A(_01064_),
    .B(_01084_),
    .C(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__a21o_1 _07028_ (.A1(net1525),
    .A2(net153),
    .B1(_01090_),
    .X(_01096_));
 sky130_fd_sc_hd__nand3_1 _07029_ (.A(net1525),
    .B(net153),
    .C(_01090_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(_01096_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _07031_ (.A(net1456),
    .B(net1913),
    .Y(_01099_));
 sky130_fd_sc_hd__xor2_1 _07032_ (.A(_01098_),
    .B(_01099_),
    .X(_01100_));
 sky130_fd_sc_hd__a21o_1 _07033_ (.A1(_01064_),
    .A2(_01084_),
    .B1(_01094_),
    .X(_01101_));
 sky130_fd_sc_hd__and3_1 _07034_ (.A(_01095_),
    .B(_01100_),
    .C(_01101_),
    .X(_01102_));
 sky130_fd_sc_hd__a31o_1 _07035_ (.A1(_01064_),
    .A2(_01084_),
    .A3(_01094_),
    .B1(_01102_),
    .X(_01103_));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(_01083_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__o21ai_1 _07037_ (.A1(_01098_),
    .A2(_01099_),
    .B1(_01097_),
    .Y(_01105_));
 sky130_fd_sc_hd__xor2_1 _07038_ (.A(_01083_),
    .B(_01103_),
    .X(_01106_));
 sky130_fd_sc_hd__a21bo_1 _07039_ (.A1(_01105_),
    .A2(_01106_),
    .B1_N(_01104_),
    .X(_01107_));
 sky130_fd_sc_hd__and2b_1 _07040_ (.A_N(_01082_),
    .B(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__xnor2_2 _07041_ (.A(_01082_),
    .B(_01107_),
    .Y(_01109_));
 sky130_fd_sc_hd__xnor2_1 _07042_ (.A(_01105_),
    .B(_01106_),
    .Y(_01110_));
 sky130_fd_sc_hd__a21oi_1 _07043_ (.A1(_01095_),
    .A2(_01101_),
    .B1(_01100_),
    .Y(_01111_));
 sky130_fd_sc_hd__a21o_1 _07044_ (.A1(_01088_),
    .A2(_01092_),
    .B1(_01091_),
    .X(_01112_));
 sky130_fd_sc_hd__a22o_1 _07045_ (.A1(net929),
    .A2(net926),
    .B1(net998),
    .B2(net800),
    .X(_01113_));
 sky130_fd_sc_hd__and4_1 _07046_ (.A(net800),
    .B(net929),
    .C(net926),
    .D(net2068),
    .X(_01114_));
 sky130_fd_sc_hd__nand4_1 _07047_ (.A(net800),
    .B(net929),
    .C(net926),
    .D(net998),
    .Y(_01115_));
 sky130_fd_sc_hd__a22o_1 _07048_ (.A1(net88),
    .A2(net2349),
    .B1(net842),
    .B2(net911),
    .X(_01116_));
 sky130_fd_sc_hd__and4_1 _07049_ (.A(_01087_),
    .B(_01113_),
    .C(_01115_),
    .D(_01116_),
    .X(_01117_));
 sky130_fd_sc_hd__nand4_1 _07050_ (.A(_01087_),
    .B(_01113_),
    .C(_01115_),
    .D(_01116_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand3_2 _07051_ (.A(_01093_),
    .B(_01112_),
    .C(_01117_),
    .Y(_01119_));
 sky130_fd_sc_hd__a21oi_1 _07052_ (.A1(net776),
    .A2(net153),
    .B1(_01114_),
    .Y(_01120_));
 sky130_fd_sc_hd__and3_1 _07053_ (.A(net776),
    .B(net153),
    .C(_01114_),
    .X(_01121_));
 sky130_fd_sc_hd__nor2_1 _07054_ (.A(_01120_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__a21oi_1 _07055_ (.A1(net697),
    .A2(net1913),
    .B1(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__and3_1 _07056_ (.A(net697),
    .B(net1913),
    .C(_01122_),
    .X(_01124_));
 sky130_fd_sc_hd__nor2_1 _07057_ (.A(_01123_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__a21o_1 _07058_ (.A1(_01093_),
    .A2(_01112_),
    .B1(_01117_),
    .X(_01126_));
 sky130_fd_sc_hd__nand3_2 _07059_ (.A(_01119_),
    .B(_01125_),
    .C(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__a211o_1 _07060_ (.A1(_01119_),
    .A2(_01127_),
    .B1(_01102_),
    .C1(_01111_),
    .X(_01128_));
 sky130_fd_sc_hd__o211ai_2 _07061_ (.A1(_01102_),
    .A2(_01111_),
    .B1(_01119_),
    .C1(_01127_),
    .Y(_01129_));
 sky130_fd_sc_hd__o211ai_2 _07062_ (.A1(_01121_),
    .A2(_01124_),
    .B1(_01128_),
    .C1(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(_01128_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__and2b_1 _07064_ (.A_N(_01110_),
    .B(_01131_),
    .X(_01132_));
 sky130_fd_sc_hd__xnor2_1 _07065_ (.A(_01110_),
    .B(_01131_),
    .Y(_01133_));
 sky130_fd_sc_hd__a211o_1 _07066_ (.A1(_01128_),
    .A2(_01129_),
    .B1(_01121_),
    .C1(_01124_),
    .X(_01134_));
 sky130_fd_sc_hd__a21o_1 _07067_ (.A1(_01119_),
    .A2(_01126_),
    .B1(_01125_),
    .X(_01135_));
 sky130_fd_sc_hd__a22o_1 _07068_ (.A1(_01113_),
    .A2(_01115_),
    .B1(_01116_),
    .B2(_01087_),
    .X(_01136_));
 sky130_fd_sc_hd__nand2_1 _07069_ (.A(_01118_),
    .B(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__and4_1 _07070_ (.A(net929),
    .B(net911),
    .C(net926),
    .D(net998),
    .X(_01138_));
 sky130_fd_sc_hd__inv_2 _07071_ (.A(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__a22o_1 _07072_ (.A1(net911),
    .A2(net2337),
    .B1(net998),
    .B2(net929),
    .X(_01140_));
 sky130_fd_sc_hd__and4_1 _07073_ (.A(net88),
    .B(net842),
    .C(_01139_),
    .D(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__a21o_1 _07074_ (.A1(net833),
    .A2(net153),
    .B1(_01138_),
    .X(_01142_));
 sky130_fd_sc_hd__nand3_1 _07075_ (.A(net833),
    .B(net153),
    .C(_01138_),
    .Y(_01143_));
 sky130_fd_sc_hd__and4_1 _07076_ (.A(net776),
    .B(net1913),
    .C(_01142_),
    .D(_01143_),
    .X(_01144_));
 sky130_fd_sc_hd__a22oi_1 _07077_ (.A1(net2829),
    .A2(net1913),
    .B1(_01142_),
    .B2(_01143_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _07078_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__xnor2_1 _07079_ (.A(_01137_),
    .B(_01141_),
    .Y(_01147_));
 sky130_fd_sc_hd__a32o_1 _07080_ (.A1(_01118_),
    .A2(_01136_),
    .A3(_01141_),
    .B1(_01146_),
    .B2(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__nand3_1 _07081_ (.A(_01127_),
    .B(_01135_),
    .C(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__a31o_1 _07082_ (.A1(net833),
    .A2(net153),
    .A3(_01138_),
    .B1(_01144_),
    .X(_01150_));
 sky130_fd_sc_hd__a21o_1 _07083_ (.A1(_01127_),
    .A2(_01135_),
    .B1(_01148_),
    .X(_01151_));
 sky130_fd_sc_hd__and3_1 _07084_ (.A(_01149_),
    .B(_01150_),
    .C(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__a21bo_1 _07085_ (.A1(_01150_),
    .A2(_01151_),
    .B1_N(_01149_),
    .X(_01153_));
 sky130_fd_sc_hd__a21oi_1 _07086_ (.A1(_01130_),
    .A2(_01134_),
    .B1(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__a21o_1 _07087_ (.A1(_01130_),
    .A2(_01134_),
    .B1(_01153_),
    .X(_01155_));
 sky130_fd_sc_hd__and3_1 _07088_ (.A(_01130_),
    .B(_01134_),
    .C(_01153_),
    .X(_01156_));
 sky130_fd_sc_hd__a21oi_1 _07089_ (.A1(_01149_),
    .A2(_01151_),
    .B1(_01150_),
    .Y(_01157_));
 sky130_fd_sc_hd__a22oi_1 _07090_ (.A1(net88),
    .A2(net842),
    .B1(_01139_),
    .B2(_01140_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _07091_ (.A(_01141_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__and4_1 _07092_ (.A(net911),
    .B(net88),
    .C(net2337),
    .D(net998),
    .X(_01160_));
 sky130_fd_sc_hd__a21oi_1 _07093_ (.A1(net800),
    .A2(net153),
    .B1(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__and3_1 _07094_ (.A(net800),
    .B(net153),
    .C(_01160_),
    .X(_01162_));
 sky130_fd_sc_hd__or2_1 _07095_ (.A(_01161_),
    .B(_01162_),
    .X(_01163_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(net2266),
    .B(net1913),
    .Y(_01164_));
 sky130_fd_sc_hd__xor2_1 _07097_ (.A(_01163_),
    .B(_01164_),
    .X(_01165_));
 sky130_fd_sc_hd__nand2_1 _07098_ (.A(_01159_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__xnor2_1 _07099_ (.A(_01146_),
    .B(_01147_),
    .Y(_01167_));
 sky130_fd_sc_hd__o21bai_1 _07100_ (.A1(_01161_),
    .A2(_01164_),
    .B1_N(_01162_),
    .Y(_01168_));
 sky130_fd_sc_hd__xor2_1 _07101_ (.A(_01166_),
    .B(_01167_),
    .X(_01169_));
 sky130_fd_sc_hd__and2_1 _07102_ (.A(_01168_),
    .B(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__o21bai_1 _07103_ (.A1(_01166_),
    .A2(_01167_),
    .B1_N(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__nor3b_1 _07104_ (.A(_01152_),
    .B(_01157_),
    .C_N(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__o21bai_2 _07105_ (.A1(_01152_),
    .A2(_01157_),
    .B1_N(_01171_),
    .Y(_01173_));
 sky130_fd_sc_hd__inv_2 _07106_ (.A(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _07107_ (.A(_01168_),
    .B(_01169_),
    .Y(_01175_));
 sky130_fd_sc_hd__or2_1 _07108_ (.A(_01170_),
    .B(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__xor2_1 _07109_ (.A(_01159_),
    .B(_01165_),
    .X(_01177_));
 sky130_fd_sc_hd__and4_1 _07110_ (.A(net2291),
    .B(net929),
    .C(net153),
    .D(net1913),
    .X(_01178_));
 sky130_fd_sc_hd__a22oi_1 _07111_ (.A1(net88),
    .A2(net2337),
    .B1(net998),
    .B2(net911),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _07112_ (.A(_01160_),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__a22o_1 _07113_ (.A1(net2168),
    .A2(net153),
    .B1(net1913),
    .B2(net2291),
    .X(_01181_));
 sky130_fd_sc_hd__and2b_1 _07114_ (.A_N(_01178_),
    .B(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__a21o_1 _07115_ (.A1(_01180_),
    .A2(_01181_),
    .B1(_01178_),
    .X(_01183_));
 sky130_fd_sc_hd__xnor2_1 _07116_ (.A(_01177_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__xnor2_1 _07117_ (.A(_01180_),
    .B(_01182_),
    .Y(_01185_));
 sky130_fd_sc_hd__and4_1 _07118_ (.A(net2168),
    .B(net911),
    .C(net153),
    .D(net1913),
    .X(_01186_));
 sky130_fd_sc_hd__inv_2 _07119_ (.A(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__a22o_1 _07120_ (.A1(net2136),
    .A2(net153),
    .B1(net1913),
    .B2(net2168),
    .X(_01188_));
 sky130_fd_sc_hd__and4b_1 _07121_ (.A_N(_01186_),
    .B(_01188_),
    .C(net88),
    .D(net998),
    .X(_01189_));
 sky130_fd_sc_hd__nor2_1 _07122_ (.A(_01186_),
    .B(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _07123_ (.A(_01185_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__a22oi_1 _07124_ (.A1(net88),
    .A2(net2066),
    .B1(_01187_),
    .B2(_01188_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _07125_ (.A(_01189_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__and4_1 _07126_ (.A(net911),
    .B(net88),
    .C(net153),
    .D(net1913),
    .X(_01194_));
 sky130_fd_sc_hd__and2_1 _07127_ (.A(_01193_),
    .B(_01194_),
    .X(_01195_));
 sky130_fd_sc_hd__xnor2_1 _07128_ (.A(_01185_),
    .B(_01190_),
    .Y(_01196_));
 sky130_fd_sc_hd__inv_2 _07129_ (.A(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__a21oi_1 _07130_ (.A1(_01195_),
    .A2(_01197_),
    .B1(_01191_),
    .Y(_01198_));
 sky130_fd_sc_hd__or2_1 _07131_ (.A(_01184_),
    .B(_01198_),
    .X(_01199_));
 sky130_fd_sc_hd__a21boi_1 _07132_ (.A1(_01177_),
    .A2(_01183_),
    .B1_N(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _07133_ (.A(_01176_),
    .B(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__or2_1 _07134_ (.A(_01176_),
    .B(_01200_),
    .X(_01202_));
 sky130_fd_sc_hd__or3_1 _07135_ (.A(_01172_),
    .B(_01174_),
    .C(_01202_),
    .X(_01203_));
 sky130_fd_sc_hd__a21oi_1 _07136_ (.A1(_01173_),
    .A2(_01201_),
    .B1(_01172_),
    .Y(_01204_));
 sky130_fd_sc_hd__a211o_1 _07137_ (.A1(_01173_),
    .A2(_01201_),
    .B1(_01156_),
    .C1(_01172_),
    .X(_01205_));
 sky130_fd_sc_hd__and3_1 _07138_ (.A(_01133_),
    .B(_01155_),
    .C(_01205_),
    .X(_01206_));
 sky130_fd_sc_hd__a31o_1 _07139_ (.A1(_01133_),
    .A2(_01155_),
    .A3(_01205_),
    .B1(_01132_),
    .X(_01207_));
 sky130_fd_sc_hd__a21o_1 _07140_ (.A1(_01109_),
    .A2(_01207_),
    .B1(_01108_),
    .X(_01208_));
 sky130_fd_sc_hd__a31o_1 _07141_ (.A1(_01080_),
    .A2(_01081_),
    .A3(_01208_),
    .B1(_01079_),
    .X(_01209_));
 sky130_fd_sc_hd__xor2_2 _07142_ (.A(_01023_),
    .B(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(net725),
    .B(net779),
    .Y(_01211_));
 sky130_fd_sc_hd__a22o_1 _07144_ (.A1(net920),
    .A2(net1853),
    .B1(net779),
    .B2(net725),
    .X(_01212_));
 sky130_fd_sc_hd__and3_1 _07145_ (.A(net725),
    .B(net1853),
    .C(net779),
    .X(_01213_));
 sky130_fd_sc_hd__a21bo_1 _07146_ (.A1(net920),
    .A2(_01213_),
    .B1_N(_01212_),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_1 _07147_ (.A(net1504),
    .B(net2114),
    .Y(_01215_));
 sky130_fd_sc_hd__xnor2_1 _07148_ (.A(_01214_),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__and4_1 _07149_ (.A(net920),
    .B(net2272),
    .C(net1853),
    .D(net779),
    .X(_01217_));
 sky130_fd_sc_hd__a22o_1 _07150_ (.A1(net2272),
    .A2(net1853),
    .B1(net779),
    .B2(net920),
    .X(_01218_));
 sky130_fd_sc_hd__inv_2 _07151_ (.A(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__and4b_1 _07152_ (.A_N(_01217_),
    .B(_01218_),
    .C(net725),
    .D(net2114),
    .X(_01220_));
 sky130_fd_sc_hd__nor2_1 _07153_ (.A(_01217_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__or2_1 _07154_ (.A(_01216_),
    .B(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__xnor2_1 _07155_ (.A(_01216_),
    .B(_01221_),
    .Y(_01223_));
 sky130_fd_sc_hd__o2bb2a_1 _07156_ (.A1_N(net725),
    .A2_N(net2114),
    .B1(_01217_),
    .B2(_01219_),
    .X(_01224_));
 sky130_fd_sc_hd__or2_1 _07157_ (.A(_01220_),
    .B(_01224_),
    .X(_01225_));
 sky130_fd_sc_hd__nand4_1 _07158_ (.A(net2272),
    .B(net2110),
    .C(net1853),
    .D(net2219),
    .Y(_01226_));
 sky130_fd_sc_hd__a22o_1 _07159_ (.A1(net2110),
    .A2(net1853),
    .B1(net2219),
    .B2(net2272),
    .X(_01227_));
 sky130_fd_sc_hd__nand2_1 _07160_ (.A(_01226_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(net920),
    .B(net2114),
    .Y(_01229_));
 sky130_fd_sc_hd__o21ai_1 _07162_ (.A1(_01228_),
    .A2(_01229_),
    .B1(_01226_),
    .Y(_01230_));
 sky130_fd_sc_hd__and2b_1 _07163_ (.A_N(_01225_),
    .B(_01230_),
    .X(_01231_));
 sky130_fd_sc_hd__and2b_1 _07164_ (.A_N(_01230_),
    .B(_01225_),
    .X(_01232_));
 sky130_fd_sc_hd__nor2_1 _07165_ (.A(_01231_),
    .B(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(net1504),
    .B(net145),
    .Y(_01234_));
 sky130_fd_sc_hd__a31oi_1 _07167_ (.A1(net1504),
    .A2(net145),
    .A3(_01233_),
    .B1(_01231_),
    .Y(_01235_));
 sky130_fd_sc_hd__or2_1 _07168_ (.A(_01223_),
    .B(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(_01223_),
    .B(_01235_),
    .Y(_01237_));
 sky130_fd_sc_hd__and2_1 _07170_ (.A(_01236_),
    .B(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__xnor2_2 _07171_ (.A(_01233_),
    .B(_01234_),
    .Y(_01239_));
 sky130_fd_sc_hd__xnor2_1 _07172_ (.A(_01228_),
    .B(_01229_),
    .Y(_01240_));
 sky130_fd_sc_hd__and4_1 _07173_ (.A(net2110),
    .B(net962),
    .C(net1853),
    .D(net779),
    .X(_01241_));
 sky130_fd_sc_hd__a22o_1 _07174_ (.A1(net962),
    .A2(net1853),
    .B1(net779),
    .B2(net2110),
    .X(_01242_));
 sky130_fd_sc_hd__nand2b_1 _07175_ (.A_N(_01241_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _07176_ (.A(net2272),
    .B(net2114),
    .Y(_01244_));
 sky130_fd_sc_hd__a31o_1 _07177_ (.A1(net2272),
    .A2(net2114),
    .A3(_01242_),
    .B1(_01241_),
    .X(_01245_));
 sky130_fd_sc_hd__nand2b_1 _07178_ (.A_N(_01240_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hd__xor2_1 _07179_ (.A(_01240_),
    .B(_01245_),
    .X(_01247_));
 sky130_fd_sc_hd__a22oi_2 _07180_ (.A1(net725),
    .A2(net145),
    .B1(net824),
    .B2(net1504),
    .Y(_01248_));
 sky130_fd_sc_hd__and4_2 _07181_ (.A(net1504),
    .B(net725),
    .C(net145),
    .D(net824),
    .X(_01249_));
 sky130_fd_sc_hd__nor2_1 _07182_ (.A(_01248_),
    .B(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__o31a_1 _07183_ (.A1(_01247_),
    .A2(_01248_),
    .A3(_01249_),
    .B1(_01246_),
    .X(_01251_));
 sky130_fd_sc_hd__and2b_1 _07184_ (.A_N(_01251_),
    .B(_01239_),
    .X(_01252_));
 sky130_fd_sc_hd__xnor2_2 _07185_ (.A(_01239_),
    .B(_01251_),
    .Y(_01253_));
 sky130_fd_sc_hd__a21oi_1 _07186_ (.A1(_01249_),
    .A2(_01253_),
    .B1(_01252_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2b_1 _07187_ (.A_N(_01254_),
    .B(_01238_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2b_1 _07188_ (.A_N(_01238_),
    .B(_01254_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_01255_),
    .B(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__xnor2_2 _07190_ (.A(_01249_),
    .B(_01253_),
    .Y(_01258_));
 sky130_fd_sc_hd__xnor2_1 _07191_ (.A(_01247_),
    .B(_01250_),
    .Y(_01259_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(_01243_),
    .B(_01244_),
    .Y(_01260_));
 sky130_fd_sc_hd__and4_1 _07193_ (.A(net962),
    .B(net887),
    .C(net1853),
    .D(net779),
    .X(_01261_));
 sky130_fd_sc_hd__a22o_1 _07194_ (.A1(net887),
    .A2(net1853),
    .B1(net779),
    .B2(net962),
    .X(_01262_));
 sky130_fd_sc_hd__nand2b_1 _07195_ (.A_N(_01261_),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(net2110),
    .B(net2114),
    .Y(_01264_));
 sky130_fd_sc_hd__a31o_1 _07197_ (.A1(net2110),
    .A2(net2114),
    .A3(_01262_),
    .B1(_01261_),
    .X(_01265_));
 sky130_fd_sc_hd__and2b_1 _07198_ (.A_N(_01260_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__xor2_1 _07199_ (.A(_01260_),
    .B(_01265_),
    .X(_01267_));
 sky130_fd_sc_hd__a22o_1 _07200_ (.A1(net920),
    .A2(net145),
    .B1(net824),
    .B2(net725),
    .X(_01268_));
 sky130_fd_sc_hd__and4_1 _07201_ (.A(net725),
    .B(net920),
    .C(net145),
    .D(net824),
    .X(_01269_));
 sky130_fd_sc_hd__nand4_1 _07202_ (.A(net725),
    .B(net920),
    .C(net145),
    .D(net824),
    .Y(_01270_));
 sky130_fd_sc_hd__a22oi_1 _07203_ (.A1(net1504),
    .A2(net1733),
    .B1(_01268_),
    .B2(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__and4_1 _07204_ (.A(net1504),
    .B(net1733),
    .C(_01268_),
    .D(_01270_),
    .X(_01272_));
 sky130_fd_sc_hd__or2_1 _07205_ (.A(_01271_),
    .B(_01272_),
    .X(_01273_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_01267_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__o21ai_2 _07207_ (.A1(_01266_),
    .A2(_01274_),
    .B1(_01259_),
    .Y(_01275_));
 sky130_fd_sc_hd__or3_2 _07208_ (.A(_01259_),
    .B(_01266_),
    .C(_01274_),
    .X(_01276_));
 sky130_fd_sc_hd__o211ai_4 _07209_ (.A1(_01269_),
    .A2(_01272_),
    .B1(_01275_),
    .C1(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _07210_ (.A(_01275_),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2b_1 _07211_ (.A_N(_01258_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _07212_ (.A(_01257_),
    .B(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__and2_1 _07213_ (.A(_01257_),
    .B(_01279_),
    .X(_01281_));
 sky130_fd_sc_hd__or2_1 _07214_ (.A(_01280_),
    .B(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__a211o_1 _07215_ (.A1(_01275_),
    .A2(_01276_),
    .B1(_01269_),
    .C1(_01272_),
    .X(_01283_));
 sky130_fd_sc_hd__xor2_1 _07216_ (.A(_01267_),
    .B(_01273_),
    .X(_01284_));
 sky130_fd_sc_hd__xnor2_2 _07217_ (.A(_01263_),
    .B(_01264_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand4_2 _07218_ (.A(net887),
    .B(net81),
    .C(net1853),
    .D(net779),
    .Y(_01286_));
 sky130_fd_sc_hd__a22o_1 _07219_ (.A1(net81),
    .A2(net1853),
    .B1(net779),
    .B2(net887),
    .X(_01287_));
 sky130_fd_sc_hd__nand4_2 _07220_ (.A(net962),
    .B(net2114),
    .C(_01286_),
    .D(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(_01286_),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__and2b_1 _07222_ (.A_N(_01285_),
    .B(_01289_),
    .X(_01290_));
 sky130_fd_sc_hd__xor2_2 _07223_ (.A(_01285_),
    .B(_01289_),
    .X(_01291_));
 sky130_fd_sc_hd__a22o_1 _07224_ (.A1(net2272),
    .A2(net145),
    .B1(net824),
    .B2(net920),
    .X(_01292_));
 sky130_fd_sc_hd__nand4_2 _07225_ (.A(net920),
    .B(net2272),
    .C(net145),
    .D(net824),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_2 _07226_ (.A(_01292_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(net725),
    .B(net1733),
    .Y(_01295_));
 sky130_fd_sc_hd__xnor2_2 _07228_ (.A(_01294_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _07229_ (.A(_01291_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21a_1 _07230_ (.A1(_01290_),
    .A2(_01297_),
    .B1(_01284_),
    .X(_01298_));
 sky130_fd_sc_hd__or3_1 _07231_ (.A(_01284_),
    .B(_01290_),
    .C(_01297_),
    .X(_01299_));
 sky130_fd_sc_hd__nand2b_1 _07232_ (.A_N(_01298_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__o21ai_2 _07233_ (.A1(_01294_),
    .A2(_01295_),
    .B1(_01293_),
    .Y(_01301_));
 sky130_fd_sc_hd__and2b_1 _07234_ (.A_N(_01300_),
    .B(_01301_),
    .X(_01302_));
 sky130_fd_sc_hd__o211ai_4 _07235_ (.A1(_01298_),
    .A2(_01302_),
    .B1(_01277_),
    .C1(_01283_),
    .Y(_01303_));
 sky130_fd_sc_hd__xor2_2 _07236_ (.A(_01258_),
    .B(_01278_),
    .X(_01304_));
 sky130_fd_sc_hd__a211o_1 _07237_ (.A1(_01277_),
    .A2(_01283_),
    .B1(_01298_),
    .C1(_01302_),
    .X(_01305_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(_01303_),
    .B(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__xnor2_2 _07239_ (.A(_01300_),
    .B(_01301_),
    .Y(_01307_));
 sky130_fd_sc_hd__xor2_2 _07240_ (.A(_01291_),
    .B(_01296_),
    .X(_01308_));
 sky130_fd_sc_hd__a22o_1 _07241_ (.A1(net962),
    .A2(net2114),
    .B1(_01286_),
    .B2(_01287_),
    .X(_01309_));
 sky130_fd_sc_hd__and4_1 _07242_ (.A(net887),
    .B(net81),
    .C(net779),
    .D(net2114),
    .X(_01310_));
 sky130_fd_sc_hd__nand3_1 _07243_ (.A(_01288_),
    .B(_01309_),
    .C(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__a22oi_1 _07244_ (.A1(net2110),
    .A2(net145),
    .B1(net2229),
    .B2(net2272),
    .Y(_01312_));
 sky130_fd_sc_hd__and4_1 _07245_ (.A(net2272),
    .B(net2110),
    .C(net145),
    .D(net2229),
    .X(_01313_));
 sky130_fd_sc_hd__nor2_1 _07246_ (.A(_01312_),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _07247_ (.A(net920),
    .B(net1733),
    .Y(_01315_));
 sky130_fd_sc_hd__and3_1 _07248_ (.A(net920),
    .B(net1733),
    .C(_01314_),
    .X(_01316_));
 sky130_fd_sc_hd__xnor2_2 _07249_ (.A(_01314_),
    .B(_01315_),
    .Y(_01317_));
 sky130_fd_sc_hd__a21o_1 _07250_ (.A1(_01288_),
    .A2(_01309_),
    .B1(_01310_),
    .X(_01318_));
 sky130_fd_sc_hd__and3_1 _07251_ (.A(_01311_),
    .B(_01317_),
    .C(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__a21boi_2 _07252_ (.A1(_01317_),
    .A2(_01318_),
    .B1_N(_01311_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2b_1 _07253_ (.A_N(_01320_),
    .B(_01308_),
    .Y(_01321_));
 sky130_fd_sc_hd__xor2_2 _07254_ (.A(_01308_),
    .B(_01320_),
    .X(_01322_));
 sky130_fd_sc_hd__o211a_1 _07255_ (.A1(_01313_),
    .A2(_01316_),
    .B1(net1504),
    .C1(net1950),
    .X(_01323_));
 sky130_fd_sc_hd__a211oi_1 _07256_ (.A1(net1504),
    .A2(net1950),
    .B1(_01313_),
    .C1(_01316_),
    .Y(_01324_));
 sky130_fd_sc_hd__or2_1 _07257_ (.A(_01323_),
    .B(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__o21ai_2 _07258_ (.A1(_01322_),
    .A2(_01325_),
    .B1(_01321_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _07259_ (.A(_01307_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__xor2_2 _07260_ (.A(_01307_),
    .B(_01326_),
    .X(_01328_));
 sky130_fd_sc_hd__a21bo_1 _07261_ (.A1(_01323_),
    .A2(_01328_),
    .B1_N(_01327_),
    .X(_01329_));
 sky130_fd_sc_hd__nand2b_1 _07262_ (.A_N(_01306_),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__xnor2_2 _07263_ (.A(_01306_),
    .B(_01329_),
    .Y(_01331_));
 sky130_fd_sc_hd__xnor2_2 _07264_ (.A(_01323_),
    .B(_01328_),
    .Y(_01332_));
 sky130_fd_sc_hd__xnor2_1 _07265_ (.A(_01322_),
    .B(_01325_),
    .Y(_01333_));
 sky130_fd_sc_hd__a21oi_1 _07266_ (.A1(_01311_),
    .A2(_01318_),
    .B1(_01317_),
    .Y(_01334_));
 sky130_fd_sc_hd__a22oi_1 _07267_ (.A1(net81),
    .A2(net779),
    .B1(net2114),
    .B2(net887),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_01310_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__a22o_1 _07269_ (.A1(net962),
    .A2(net145),
    .B1(net824),
    .B2(net2110),
    .X(_01337_));
 sky130_fd_sc_hd__nand4_2 _07270_ (.A(net2110),
    .B(net962),
    .C(net145),
    .D(net824),
    .Y(_01338_));
 sky130_fd_sc_hd__and2_1 _07271_ (.A(net2272),
    .B(net1733),
    .X(_01339_));
 sky130_fd_sc_hd__a21o_1 _07272_ (.A1(_01337_),
    .A2(_01338_),
    .B1(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__nand3_1 _07273_ (.A(_01337_),
    .B(_01338_),
    .C(_01339_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand3_1 _07274_ (.A(_01336_),
    .B(_01340_),
    .C(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__or3_2 _07275_ (.A(_01319_),
    .B(_01334_),
    .C(_01342_),
    .X(_01343_));
 sky130_fd_sc_hd__a21bo_1 _07276_ (.A1(_01337_),
    .A2(_01339_),
    .B1_N(_01338_),
    .X(_01344_));
 sky130_fd_sc_hd__a21oi_1 _07277_ (.A1(net725),
    .A2(net1950),
    .B1(_01344_),
    .Y(_01345_));
 sky130_fd_sc_hd__and3_1 _07278_ (.A(net725),
    .B(net1950),
    .C(_01344_),
    .X(_01346_));
 sky130_fd_sc_hd__nor2_1 _07279_ (.A(_01345_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(net1504),
    .B(net890),
    .Y(_01348_));
 sky130_fd_sc_hd__xnor2_1 _07281_ (.A(_01347_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__o21ai_1 _07282_ (.A1(_01319_),
    .A2(_01334_),
    .B1(_01342_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand3_2 _07283_ (.A(_01343_),
    .B(_01349_),
    .C(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(_01343_),
    .B(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2b_1 _07285_ (.A_N(_01333_),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__xnor2_1 _07286_ (.A(_01333_),
    .B(_01352_),
    .Y(_01354_));
 sky130_fd_sc_hd__a31o_1 _07287_ (.A1(net1504),
    .A2(net890),
    .A3(_01347_),
    .B1(_01346_),
    .X(_01355_));
 sky130_fd_sc_hd__a21bo_1 _07288_ (.A1(_01354_),
    .A2(_01355_),
    .B1_N(_01353_),
    .X(_01356_));
 sky130_fd_sc_hd__and2b_1 _07289_ (.A_N(_01332_),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__xnor2_2 _07290_ (.A(_01332_),
    .B(_01356_),
    .Y(_01358_));
 sky130_fd_sc_hd__xnor2_1 _07291_ (.A(_01354_),
    .B(_01355_),
    .Y(_01359_));
 sky130_fd_sc_hd__a21o_1 _07292_ (.A1(_01343_),
    .A2(_01350_),
    .B1(_01349_),
    .X(_01360_));
 sky130_fd_sc_hd__a21o_1 _07293_ (.A1(_01340_),
    .A2(_01341_),
    .B1(_01336_),
    .X(_01361_));
 sky130_fd_sc_hd__a22o_1 _07294_ (.A1(net887),
    .A2(net145),
    .B1(net824),
    .B2(net962),
    .X(_01362_));
 sky130_fd_sc_hd__nand4_1 _07295_ (.A(net962),
    .B(net887),
    .C(net145),
    .D(net824),
    .Y(_01363_));
 sky130_fd_sc_hd__and2_1 _07296_ (.A(net2110),
    .B(net1733),
    .X(_01364_));
 sky130_fd_sc_hd__a21oi_1 _07297_ (.A1(_01362_),
    .A2(_01363_),
    .B1(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__and3_1 _07298_ (.A(_01362_),
    .B(_01363_),
    .C(_01364_),
    .X(_01366_));
 sky130_fd_sc_hd__and4bb_1 _07299_ (.A_N(_01365_),
    .B_N(_01366_),
    .C(net81),
    .D(net2114),
    .X(_01367_));
 sky130_fd_sc_hd__nand3_1 _07300_ (.A(_01342_),
    .B(_01361_),
    .C(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__a21bo_1 _07301_ (.A1(_01362_),
    .A2(_01364_),
    .B1_N(_01363_),
    .X(_01369_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(net920),
    .B(net1950),
    .Y(_01370_));
 sky130_fd_sc_hd__and3_1 _07303_ (.A(net920),
    .B(net1950),
    .C(_01369_),
    .X(_01371_));
 sky130_fd_sc_hd__xnor2_1 _07304_ (.A(_01369_),
    .B(_01370_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _07305_ (.A(net1558),
    .B(net890),
    .Y(_01373_));
 sky130_fd_sc_hd__xnor2_1 _07306_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__a21o_1 _07307_ (.A1(_01342_),
    .A2(_01361_),
    .B1(_01367_),
    .X(_01375_));
 sky130_fd_sc_hd__nand3_1 _07308_ (.A(_01368_),
    .B(_01374_),
    .C(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _07309_ (.A(_01368_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand3_1 _07310_ (.A(_01351_),
    .B(_01360_),
    .C(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__a31o_1 _07311_ (.A1(net3699),
    .A2(net890),
    .A3(_01372_),
    .B1(_01371_),
    .X(_01379_));
 sky130_fd_sc_hd__a21o_1 _07312_ (.A1(_01351_),
    .A2(_01360_),
    .B1(_01377_),
    .X(_01380_));
 sky130_fd_sc_hd__and3_1 _07313_ (.A(_01378_),
    .B(_01379_),
    .C(_01380_),
    .X(_01381_));
 sky130_fd_sc_hd__a31o_1 _07314_ (.A1(_01351_),
    .A2(_01360_),
    .A3(_01377_),
    .B1(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__and2b_1 _07315_ (.A_N(_01359_),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__xnor2_1 _07316_ (.A(_01359_),
    .B(_01382_),
    .Y(_01384_));
 sky130_fd_sc_hd__a21oi_1 _07317_ (.A1(_01378_),
    .A2(_01380_),
    .B1(_01379_),
    .Y(_01385_));
 sky130_fd_sc_hd__a21o_1 _07318_ (.A1(_01368_),
    .A2(_01375_),
    .B1(_01374_),
    .X(_01386_));
 sky130_fd_sc_hd__o2bb2a_1 _07319_ (.A1_N(net81),
    .A2_N(net2114),
    .B1(_01365_),
    .B2(_01366_),
    .X(_01387_));
 sky130_fd_sc_hd__nor2_1 _07320_ (.A(_01367_),
    .B(_01387_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand2_1 _07321_ (.A(net2469),
    .B(net890),
    .Y(_01389_));
 sky130_fd_sc_hd__and3_1 _07322_ (.A(net887),
    .B(net81),
    .C(net824),
    .X(_01390_));
 sky130_fd_sc_hd__nand2_1 _07323_ (.A(net962),
    .B(net1733),
    .Y(_01391_));
 sky130_fd_sc_hd__a22o_1 _07324_ (.A1(net81),
    .A2(net145),
    .B1(net824),
    .B2(net2060),
    .X(_01392_));
 sky130_fd_sc_hd__a21bo_1 _07325_ (.A1(net1369),
    .A2(_01390_),
    .B1_N(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__a32o_1 _07326_ (.A1(net962),
    .A2(net1733),
    .A3(_01392_),
    .B1(_01390_),
    .B2(net1369),
    .X(_01394_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(net2272),
    .B(net1950),
    .Y(_01395_));
 sky130_fd_sc_hd__and3_1 _07328_ (.A(net2272),
    .B(net1950),
    .C(_01394_),
    .X(_01396_));
 sky130_fd_sc_hd__xnor2_1 _07329_ (.A(_01394_),
    .B(_01395_),
    .Y(_01397_));
 sky130_fd_sc_hd__xnor2_1 _07330_ (.A(_01389_),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__and2_1 _07331_ (.A(_01388_),
    .B(_01398_),
    .X(_01399_));
 sky130_fd_sc_hd__and3_1 _07332_ (.A(_01376_),
    .B(_01386_),
    .C(_01399_),
    .X(_01400_));
 sky130_fd_sc_hd__nand3_1 _07333_ (.A(_01376_),
    .B(_01386_),
    .C(_01399_),
    .Y(_01401_));
 sky130_fd_sc_hd__a31oi_1 _07334_ (.A1(net2469),
    .A2(net890),
    .A3(_01397_),
    .B1(_01396_),
    .Y(_01402_));
 sky130_fd_sc_hd__a21oi_1 _07335_ (.A1(_01376_),
    .A2(_01386_),
    .B1(_01399_),
    .Y(_01403_));
 sky130_fd_sc_hd__or3_2 _07336_ (.A(_01400_),
    .B(_01402_),
    .C(_01403_),
    .X(_01404_));
 sky130_fd_sc_hd__a211oi_1 _07337_ (.A1(_01401_),
    .A2(_01404_),
    .B1(_01381_),
    .C1(_01385_),
    .Y(_01405_));
 sky130_fd_sc_hd__o211ai_1 _07338_ (.A1(_01381_),
    .A2(_01385_),
    .B1(_01401_),
    .C1(_01404_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2b_1 _07339_ (.A_N(_01405_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__o21ai_1 _07340_ (.A1(_01400_),
    .A2(_01403_),
    .B1(_01402_),
    .Y(_01408_));
 sky130_fd_sc_hd__xnor2_1 _07341_ (.A(_01388_),
    .B(_01398_),
    .Y(_01409_));
 sky130_fd_sc_hd__xor2_1 _07342_ (.A(_01391_),
    .B(_01393_),
    .X(_01410_));
 sky130_fd_sc_hd__and4_1 _07343_ (.A(net887),
    .B(net81),
    .C(net824),
    .D(net1733),
    .X(_01411_));
 sky130_fd_sc_hd__inv_2 _07344_ (.A(_01411_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _07345_ (.A(net2110),
    .B(net1950),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _07346_ (.A(_01412_),
    .B(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__xnor2_1 _07347_ (.A(_01411_),
    .B(_01413_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(net2272),
    .B(net890),
    .Y(_01416_));
 sky130_fd_sc_hd__xnor2_1 _07349_ (.A(_01415_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(_01410_),
    .B(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _07351_ (.A(_01409_),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__a31o_1 _07352_ (.A1(net2272),
    .A2(net890),
    .A3(_01415_),
    .B1(_01414_),
    .X(_01420_));
 sky130_fd_sc_hd__xor2_1 _07353_ (.A(_01409_),
    .B(_01418_),
    .X(_01421_));
 sky130_fd_sc_hd__a21o_1 _07354_ (.A1(_01420_),
    .A2(_01421_),
    .B1(_01419_),
    .X(_01422_));
 sky130_fd_sc_hd__and3_1 _07355_ (.A(_01404_),
    .B(_01408_),
    .C(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__a21o_1 _07356_ (.A1(_01404_),
    .A2(_01408_),
    .B1(_01422_),
    .X(_01424_));
 sky130_fd_sc_hd__and2b_1 _07357_ (.A_N(_01423_),
    .B(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__xnor2_1 _07358_ (.A(_01420_),
    .B(_01421_),
    .Y(_01426_));
 sky130_fd_sc_hd__or2_1 _07359_ (.A(_01410_),
    .B(_01417_),
    .X(_01427_));
 sky130_fd_sc_hd__and2_1 _07360_ (.A(_01418_),
    .B(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__and4_1 _07361_ (.A(net2110),
    .B(net962),
    .C(net1950),
    .D(net890),
    .X(_01429_));
 sky130_fd_sc_hd__inv_2 _07362_ (.A(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__a22o_1 _07363_ (.A1(net81),
    .A2(net824),
    .B1(net1733),
    .B2(net887),
    .X(_01431_));
 sky130_fd_sc_hd__a22o_1 _07364_ (.A1(net962),
    .A2(net1950),
    .B1(net890),
    .B2(net2110),
    .X(_01432_));
 sky130_fd_sc_hd__or4bb_1 _07365_ (.A(_01411_),
    .B(_01429_),
    .C_N(_01431_),
    .D_N(_01432_),
    .X(_01433_));
 sky130_fd_sc_hd__nand2_1 _07366_ (.A(_01430_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _07367_ (.A(_01428_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__xnor2_1 _07368_ (.A(_01428_),
    .B(_01434_),
    .Y(_01436_));
 sky130_fd_sc_hd__a22o_1 _07369_ (.A1(_01412_),
    .A2(_01431_),
    .B1(_01432_),
    .B2(_01430_),
    .X(_01437_));
 sky130_fd_sc_hd__and4_1 _07370_ (.A(net962),
    .B(net887),
    .C(net1950),
    .D(net890),
    .X(_01438_));
 sky130_fd_sc_hd__a22o_1 _07371_ (.A1(net887),
    .A2(net1950),
    .B1(net890),
    .B2(net2213),
    .X(_01439_));
 sky130_fd_sc_hd__inv_2 _07372_ (.A(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__and4b_1 _07373_ (.A_N(_01438_),
    .B(_01439_),
    .C(net81),
    .D(net1733),
    .X(_01441_));
 sky130_fd_sc_hd__or2_1 _07374_ (.A(_01438_),
    .B(_01441_),
    .X(_01442_));
 sky130_fd_sc_hd__and3_1 _07375_ (.A(_01433_),
    .B(_01437_),
    .C(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__o2bb2a_1 _07376_ (.A1_N(net81),
    .A2_N(net1733),
    .B1(_01438_),
    .B2(_01440_),
    .X(_01444_));
 sky130_fd_sc_hd__nor2_1 _07377_ (.A(_01441_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__and4_1 _07378_ (.A(net887),
    .B(net81),
    .C(net1950),
    .D(net2156),
    .X(_01446_));
 sky130_fd_sc_hd__and2_1 _07379_ (.A(_01445_),
    .B(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__a21oi_1 _07380_ (.A1(_01433_),
    .A2(_01437_),
    .B1(_01442_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _07381_ (.A(_01443_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__and2_1 _07382_ (.A(_01447_),
    .B(_01449_),
    .X(_01450_));
 sky130_fd_sc_hd__nor2_1 _07383_ (.A(_01443_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__o21bai_2 _07384_ (.A1(_01443_),
    .A2(_01450_),
    .B1_N(_01436_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21oi_2 _07385_ (.A1(_01435_),
    .A2(_01452_),
    .B1(_01426_),
    .Y(_01453_));
 sky130_fd_sc_hd__a21o_1 _07386_ (.A1(_01424_),
    .A2(_01453_),
    .B1(_01423_),
    .X(_01454_));
 sky130_fd_sc_hd__a21o_1 _07387_ (.A1(_01406_),
    .A2(_01454_),
    .B1(_01405_),
    .X(_01455_));
 sky130_fd_sc_hd__a21o_1 _07388_ (.A1(_01384_),
    .A2(_01455_),
    .B1(_01383_),
    .X(_01456_));
 sky130_fd_sc_hd__a21o_1 _07389_ (.A1(_01358_),
    .A2(_01456_),
    .B1(_01357_),
    .X(_01457_));
 sky130_fd_sc_hd__a21boi_2 _07390_ (.A1(_01331_),
    .A2(_01457_),
    .B1_N(_01330_),
    .Y(_01458_));
 sky130_fd_sc_hd__a21o_1 _07391_ (.A1(_01303_),
    .A2(_01458_),
    .B1(_01304_),
    .X(_01459_));
 sky130_fd_sc_hd__a211oi_1 _07392_ (.A1(_01303_),
    .A2(_01458_),
    .B1(_01304_),
    .C1(_01282_),
    .Y(_01460_));
 sky130_fd_sc_hd__xnor2_1 _07393_ (.A(_01282_),
    .B(_01459_),
    .Y(_01461_));
 sky130_fd_sc_hd__xnor2_1 _07394_ (.A(_00952_),
    .B(_01210_),
    .Y(_01462_));
 sky130_fd_sc_hd__or2_1 _07395_ (.A(_01461_),
    .B(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__a21bo_1 _07396_ (.A1(_00952_),
    .A2(_01210_),
    .B1_N(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(net482),
    .B(net140),
    .Y(_01465_));
 sky130_fd_sc_hd__a22o_1 _07398_ (.A1(net1883),
    .A2(net1777),
    .B1(net140),
    .B2(net482),
    .X(_01466_));
 sky130_fd_sc_hd__and3_1 _07399_ (.A(net1883),
    .B(net1777),
    .C(net140),
    .X(_01467_));
 sky130_fd_sc_hd__a21bo_1 _07400_ (.A1(net482),
    .A2(_01467_),
    .B1_N(_01466_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(net1411),
    .B(net1801),
    .Y(_01469_));
 sky130_fd_sc_hd__xor2_1 _07402_ (.A(_01468_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__and4_1 _07403_ (.A(net1883),
    .B(net2082),
    .C(net1777),
    .D(net140),
    .X(_01471_));
 sky130_fd_sc_hd__inv_2 _07404_ (.A(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__a22o_1 _07405_ (.A1(net2082),
    .A2(net1777),
    .B1(net140),
    .B2(net1883),
    .X(_01473_));
 sky130_fd_sc_hd__and4_1 _07406_ (.A(net482),
    .B(net1801),
    .C(_01472_),
    .D(_01473_),
    .X(_01474_));
 sky130_fd_sc_hd__o21ai_2 _07407_ (.A1(_01471_),
    .A2(_01474_),
    .B1(_01470_),
    .Y(_01475_));
 sky130_fd_sc_hd__or3_1 _07408_ (.A(_01470_),
    .B(_01471_),
    .C(_01474_),
    .X(_01476_));
 sky130_fd_sc_hd__nand2_1 _07409_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__a22oi_1 _07410_ (.A1(net482),
    .A2(net1801),
    .B1(_01472_),
    .B2(_01473_),
    .Y(_01478_));
 sky130_fd_sc_hd__or2_1 _07411_ (.A(_01474_),
    .B(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__nand4_1 _07412_ (.A(net2082),
    .B(net1974),
    .C(net1777),
    .D(net140),
    .Y(_01480_));
 sky130_fd_sc_hd__a22o_1 _07413_ (.A1(net1974),
    .A2(net1777),
    .B1(net140),
    .B2(net2082),
    .X(_01481_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_01480_),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _07415_ (.A(net1883),
    .B(net1801),
    .Y(_01483_));
 sky130_fd_sc_hd__o21ai_1 _07416_ (.A1(_01482_),
    .A2(_01483_),
    .B1(_01480_),
    .Y(_01484_));
 sky130_fd_sc_hd__and2b_1 _07417_ (.A_N(_01479_),
    .B(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__and2b_1 _07418_ (.A_N(_01484_),
    .B(_01479_),
    .X(_01486_));
 sky130_fd_sc_hd__nor2_1 _07419_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _07420_ (.A(net1411),
    .B(net1168),
    .Y(_01488_));
 sky130_fd_sc_hd__a31oi_1 _07421_ (.A1(net1411),
    .A2(net1168),
    .A3(_01487_),
    .B1(_01485_),
    .Y(_01489_));
 sky130_fd_sc_hd__or2_1 _07422_ (.A(_01477_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _07423_ (.A(_01477_),
    .B(_01489_),
    .Y(_01491_));
 sky130_fd_sc_hd__and2_1 _07424_ (.A(_01490_),
    .B(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__xnor2_1 _07425_ (.A(_01487_),
    .B(_01488_),
    .Y(_01493_));
 sky130_fd_sc_hd__xnor2_1 _07426_ (.A(_01482_),
    .B(_01483_),
    .Y(_01494_));
 sky130_fd_sc_hd__and4_1 _07427_ (.A(net1974),
    .B(net1694),
    .C(net1777),
    .D(net140),
    .X(_01495_));
 sky130_fd_sc_hd__inv_2 _07428_ (.A(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__a22o_1 _07429_ (.A1(net1694),
    .A2(net1777),
    .B1(net140),
    .B2(net1974),
    .X(_01497_));
 sky130_fd_sc_hd__and4_1 _07430_ (.A(net2082),
    .B(net1801),
    .C(_01496_),
    .D(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__or2_1 _07431_ (.A(_01495_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2b_1 _07432_ (.A_N(_01494_),
    .B(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__and2b_1 _07433_ (.A_N(_01499_),
    .B(_01494_),
    .X(_01501_));
 sky130_fd_sc_hd__or2_1 _07434_ (.A(_01500_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__a22oi_1 _07435_ (.A1(net482),
    .A2(net1168),
    .B1(net1737),
    .B2(net1411),
    .Y(_01503_));
 sky130_fd_sc_hd__and4_1 _07436_ (.A(net1411),
    .B(net482),
    .C(net1168),
    .D(net1737),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_1 _07437_ (.A(_01503_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__and2b_1 _07438_ (.A_N(_01502_),
    .B(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_01500_),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__o21a_1 _07440_ (.A1(_01500_),
    .A2(_01506_),
    .B1(_01493_),
    .X(_01508_));
 sky130_fd_sc_hd__xnor2_1 _07441_ (.A(_01493_),
    .B(_01507_),
    .Y(_01509_));
 sky130_fd_sc_hd__a21oi_1 _07442_ (.A1(_01504_),
    .A2(_01509_),
    .B1(_01508_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2b_2 _07443_ (.A_N(_01510_),
    .B(_01492_),
    .Y(_01511_));
 sky130_fd_sc_hd__a22oi_1 _07444_ (.A1(net482),
    .A2(net1777),
    .B1(net140),
    .B2(net1411),
    .Y(_01512_));
 sky130_fd_sc_hd__and4_1 _07445_ (.A(net1411),
    .B(net482),
    .C(net1777),
    .D(net140),
    .X(_01513_));
 sky130_fd_sc_hd__nor2_1 _07446_ (.A(_01512_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__a32o_1 _07447_ (.A1(net1411),
    .A2(net1801),
    .A3(_01466_),
    .B1(_01467_),
    .B2(net482),
    .X(_01515_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(_01514_),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__or2_1 _07449_ (.A(_01514_),
    .B(_01515_),
    .X(_01517_));
 sky130_fd_sc_hd__nand2_2 _07450_ (.A(_01516_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_01475_),
    .B(_01490_),
    .Y(_01519_));
 sky130_fd_sc_hd__xnor2_2 _07452_ (.A(_01518_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand2b_1 _07453_ (.A_N(_01511_),
    .B(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__xnor2_2 _07454_ (.A(_01511_),
    .B(_01520_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2b_1 _07455_ (.A_N(_01492_),
    .B(_01510_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _07456_ (.A(_01511_),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__xnor2_1 _07457_ (.A(_01504_),
    .B(_01509_),
    .Y(_01525_));
 sky130_fd_sc_hd__xnor2_1 _07458_ (.A(_01502_),
    .B(_01505_),
    .Y(_01526_));
 sky130_fd_sc_hd__a22oi_1 _07459_ (.A1(net2082),
    .A2(net1801),
    .B1(_01496_),
    .B2(_01497_),
    .Y(_01527_));
 sky130_fd_sc_hd__or2_1 _07460_ (.A(_01498_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__and4_1 _07461_ (.A(net1694),
    .B(net740),
    .C(net1777),
    .D(net140),
    .X(_01529_));
 sky130_fd_sc_hd__a22o_1 _07462_ (.A1(net740),
    .A2(net1777),
    .B1(net140),
    .B2(net1694),
    .X(_01530_));
 sky130_fd_sc_hd__nand2b_1 _07463_ (.A_N(_01529_),
    .B(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand2_1 _07464_ (.A(net1974),
    .B(net1801),
    .Y(_01532_));
 sky130_fd_sc_hd__a31o_1 _07465_ (.A1(net1974),
    .A2(net1801),
    .A3(_01530_),
    .B1(_01529_),
    .X(_01533_));
 sky130_fd_sc_hd__or3b_1 _07466_ (.A(_01498_),
    .B(_01527_),
    .C_N(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__xor2_1 _07467_ (.A(_01528_),
    .B(_01533_),
    .X(_01535_));
 sky130_fd_sc_hd__a22o_1 _07468_ (.A1(net1883),
    .A2(net1168),
    .B1(net1737),
    .B2(net1465),
    .X(_01536_));
 sky130_fd_sc_hd__and4_1 _07469_ (.A(net1465),
    .B(net1883),
    .C(net1168),
    .D(net1737),
    .X(_01537_));
 sky130_fd_sc_hd__inv_2 _07470_ (.A(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__and2_1 _07471_ (.A(_01536_),
    .B(_01538_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2b_1 _07472_ (.A_N(_01535_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _07473_ (.A(_01534_),
    .B(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__xnor2_1 _07474_ (.A(_01526_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _07475_ (.A(_01538_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_1 _07476_ (.A1(_01526_),
    .A2(_01541_),
    .B1(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2b_1 _07477_ (.A_N(_01525_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__nor2_1 _07478_ (.A(_01524_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__and2_1 _07479_ (.A(_01524_),
    .B(_01545_),
    .X(_01547_));
 sky130_fd_sc_hd__nor2_1 _07480_ (.A(_01546_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__xnor2_1 _07481_ (.A(_01525_),
    .B(_01544_),
    .Y(_01549_));
 sky130_fd_sc_hd__xnor2_1 _07482_ (.A(_01538_),
    .B(_01542_),
    .Y(_01550_));
 sky130_fd_sc_hd__xnor2_1 _07483_ (.A(_01535_),
    .B(_01539_),
    .Y(_01551_));
 sky130_fd_sc_hd__xnor2_1 _07484_ (.A(_01531_),
    .B(_01532_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand4_2 _07485_ (.A(net740),
    .B(net761),
    .C(net1777),
    .D(net140),
    .Y(_01553_));
 sky130_fd_sc_hd__a22o_1 _07486_ (.A1(net761),
    .A2(net1777),
    .B1(net140),
    .B2(net740),
    .X(_01554_));
 sky130_fd_sc_hd__nand4_2 _07487_ (.A(net1694),
    .B(net1801),
    .C(_01553_),
    .D(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _07488_ (.A(_01553_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__and2b_1 _07489_ (.A_N(_01552_),
    .B(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__xor2_1 _07490_ (.A(_01552_),
    .B(_01556_),
    .X(_01558_));
 sky130_fd_sc_hd__a22o_1 _07491_ (.A1(net2082),
    .A2(net1168),
    .B1(net1737),
    .B2(net1883),
    .X(_01559_));
 sky130_fd_sc_hd__inv_2 _07492_ (.A(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__and4_1 _07493_ (.A(net1883),
    .B(net2082),
    .C(net1168),
    .D(net1737),
    .X(_01561_));
 sky130_fd_sc_hd__nor2_1 _07494_ (.A(_01560_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__and2b_1 _07495_ (.A_N(_01558_),
    .B(_01562_),
    .X(_01563_));
 sky130_fd_sc_hd__or2_1 _07496_ (.A(_01557_),
    .B(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__nand2_1 _07497_ (.A(_01551_),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__xnor2_1 _07498_ (.A(_01551_),
    .B(_01564_),
    .Y(_01566_));
 sky130_fd_sc_hd__and3_1 _07499_ (.A(net1411),
    .B(net1786),
    .C(_01561_),
    .X(_01567_));
 sky130_fd_sc_hd__inv_2 _07500_ (.A(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a21oi_1 _07501_ (.A1(net1411),
    .A2(net1786),
    .B1(_01561_),
    .Y(_01569_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(_01567_),
    .B(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__o21a_1 _07503_ (.A1(_01566_),
    .A2(_01570_),
    .B1(_01565_),
    .X(_01571_));
 sky130_fd_sc_hd__nor2_1 _07504_ (.A(_01550_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__xnor2_1 _07505_ (.A(_01550_),
    .B(_01571_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _07506_ (.A(_01568_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__o21a_1 _07507_ (.A1(_01572_),
    .A2(_01574_),
    .B1(_01549_),
    .X(_01575_));
 sky130_fd_sc_hd__nor3_1 _07508_ (.A(_01549_),
    .B(_01572_),
    .C(_01574_),
    .Y(_01576_));
 sky130_fd_sc_hd__or2_1 _07509_ (.A(_01575_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__xnor2_1 _07510_ (.A(_01567_),
    .B(_01573_),
    .Y(_01578_));
 sky130_fd_sc_hd__xor2_1 _07511_ (.A(_01566_),
    .B(_01570_),
    .X(_01579_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(_01558_),
    .B(_01562_),
    .Y(_01580_));
 sky130_fd_sc_hd__a22o_1 _07513_ (.A1(net1694),
    .A2(net1801),
    .B1(_01553_),
    .B2(_01554_),
    .X(_01581_));
 sky130_fd_sc_hd__and4_1 _07514_ (.A(net740),
    .B(net761),
    .C(net140),
    .D(net1801),
    .X(_01582_));
 sky130_fd_sc_hd__and3_1 _07515_ (.A(_01555_),
    .B(_01581_),
    .C(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__nand3_1 _07516_ (.A(_01555_),
    .B(_01581_),
    .C(_01582_),
    .Y(_01584_));
 sky130_fd_sc_hd__a21o_1 _07517_ (.A1(_01555_),
    .A2(_01581_),
    .B1(_01582_),
    .X(_01585_));
 sky130_fd_sc_hd__nand2_1 _07518_ (.A(net2082),
    .B(net1737),
    .Y(_01586_));
 sky130_fd_sc_hd__a22oi_1 _07519_ (.A1(net1974),
    .A2(net1168),
    .B1(net1118),
    .B2(net1411),
    .Y(_01587_));
 sky130_fd_sc_hd__and4_1 _07520_ (.A(net1411),
    .B(net1974),
    .C(net1168),
    .D(net1118),
    .X(_01588_));
 sky130_fd_sc_hd__nor2_1 _07521_ (.A(_01587_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__xnor2_1 _07522_ (.A(_01586_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__and3_1 _07523_ (.A(_01584_),
    .B(_01585_),
    .C(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__nor2_1 _07524_ (.A(_01583_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__and2b_1 _07525_ (.A_N(_01592_),
    .B(_01580_),
    .X(_01593_));
 sky130_fd_sc_hd__xnor2_1 _07526_ (.A(_01580_),
    .B(_01592_),
    .Y(_01594_));
 sky130_fd_sc_hd__o21bai_1 _07527_ (.A1(_01586_),
    .A2(_01587_),
    .B1_N(_01588_),
    .Y(_01595_));
 sky130_fd_sc_hd__and2_1 _07528_ (.A(net1411),
    .B(net815),
    .X(_01596_));
 sky130_fd_sc_hd__nor2_1 _07529_ (.A(_01595_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__and2_1 _07530_ (.A(_01595_),
    .B(_01596_),
    .X(_01598_));
 sky130_fd_sc_hd__nor2_1 _07531_ (.A(_01597_),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__and2_1 _07532_ (.A(net482),
    .B(net1786),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_1 _07533_ (.A(_01599_),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__and2_1 _07534_ (.A(_01599_),
    .B(_01600_),
    .X(_01602_));
 sky130_fd_sc_hd__nor2_1 _07535_ (.A(_01601_),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21oi_1 _07536_ (.A1(_01594_),
    .A2(_01603_),
    .B1(_01593_),
    .Y(_01604_));
 sky130_fd_sc_hd__and2b_1 _07537_ (.A_N(_01604_),
    .B(_01579_),
    .X(_01605_));
 sky130_fd_sc_hd__xnor2_1 _07538_ (.A(_01579_),
    .B(_01604_),
    .Y(_01606_));
 sky130_fd_sc_hd__o21a_1 _07539_ (.A1(_01598_),
    .A2(_01602_),
    .B1(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_1 _07540_ (.A(_01605_),
    .B(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2b_1 _07541_ (.A_N(_01608_),
    .B(_01578_),
    .Y(_01609_));
 sky130_fd_sc_hd__xnor2_1 _07542_ (.A(_01578_),
    .B(_01608_),
    .Y(_01610_));
 sky130_fd_sc_hd__nor3_1 _07543_ (.A(_01598_),
    .B(_01602_),
    .C(_01606_),
    .Y(_01611_));
 sky130_fd_sc_hd__xnor2_1 _07544_ (.A(_01594_),
    .B(_01603_),
    .Y(_01612_));
 sky130_fd_sc_hd__a21oi_1 _07545_ (.A1(_01584_),
    .A2(_01585_),
    .B1(_01590_),
    .Y(_01613_));
 sky130_fd_sc_hd__a22oi_1 _07546_ (.A1(net761),
    .A2(net1329),
    .B1(net1801),
    .B2(net740),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _07547_ (.A(_01582_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__a22o_1 _07548_ (.A1(net1694),
    .A2(net1168),
    .B1(net1118),
    .B2(net482),
    .X(_01616_));
 sky130_fd_sc_hd__nand4_1 _07549_ (.A(net482),
    .B(net1694),
    .C(net1168),
    .D(net1118),
    .Y(_01617_));
 sky130_fd_sc_hd__and2_1 _07550_ (.A(net1974),
    .B(net1737),
    .X(_01618_));
 sky130_fd_sc_hd__a21o_1 _07551_ (.A1(_01616_),
    .A2(_01617_),
    .B1(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__nand3_1 _07552_ (.A(_01616_),
    .B(_01617_),
    .C(_01618_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand3_1 _07553_ (.A(_01615_),
    .B(_01619_),
    .C(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__or3_2 _07554_ (.A(_01591_),
    .B(_01613_),
    .C(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__o21ai_1 _07555_ (.A1(_01591_),
    .A2(_01613_),
    .B1(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__a21bo_1 _07556_ (.A1(_01616_),
    .A2(_01618_),
    .B1_N(_01617_),
    .X(_01624_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(net482),
    .B(net815),
    .Y(_01625_));
 sky130_fd_sc_hd__and3_1 _07558_ (.A(net1467),
    .B(net815),
    .C(_01624_),
    .X(_01626_));
 sky130_fd_sc_hd__xnor2_1 _07559_ (.A(_01624_),
    .B(_01625_),
    .Y(_01627_));
 sky130_fd_sc_hd__and2_1 _07560_ (.A(net1883),
    .B(net1786),
    .X(_01628_));
 sky130_fd_sc_hd__nor2_1 _07561_ (.A(_01627_),
    .B(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__and2_1 _07562_ (.A(_01627_),
    .B(_01628_),
    .X(_01630_));
 sky130_fd_sc_hd__nor2_1 _07563_ (.A(_01629_),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand3_2 _07564_ (.A(_01622_),
    .B(_01623_),
    .C(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__a21o_2 _07565_ (.A1(_01622_),
    .A2(_01632_),
    .B1(_01612_),
    .X(_01633_));
 sky130_fd_sc_hd__nand3_2 _07566_ (.A(_01612_),
    .B(_01622_),
    .C(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__o211ai_4 _07567_ (.A1(_01626_),
    .A2(_01630_),
    .B1(_01633_),
    .C1(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__a211oi_2 _07568_ (.A1(_01633_),
    .A2(_01635_),
    .B1(_01607_),
    .C1(_01611_),
    .Y(_01636_));
 sky130_fd_sc_hd__o211a_1 _07569_ (.A1(_01607_),
    .A2(_01611_),
    .B1(_01633_),
    .C1(_01635_),
    .X(_01637_));
 sky130_fd_sc_hd__a211o_1 _07570_ (.A1(_01633_),
    .A2(_01634_),
    .B1(_01626_),
    .C1(_01630_),
    .X(_01638_));
 sky130_fd_sc_hd__a21o_1 _07571_ (.A1(_01622_),
    .A2(_01623_),
    .B1(_01631_),
    .X(_01639_));
 sky130_fd_sc_hd__a21o_1 _07572_ (.A1(_01619_),
    .A2(_01620_),
    .B1(_01615_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _07573_ (.A1(net740),
    .A2(net1168),
    .B1(net1118),
    .B2(net1883),
    .X(_01641_));
 sky130_fd_sc_hd__nand4_2 _07574_ (.A(net1883),
    .B(net1656),
    .C(net1168),
    .D(net1118),
    .Y(_01642_));
 sky130_fd_sc_hd__and2_1 _07575_ (.A(net1694),
    .B(net1737),
    .X(_01643_));
 sky130_fd_sc_hd__a21oi_1 _07576_ (.A1(_01641_),
    .A2(_01642_),
    .B1(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__and3_1 _07577_ (.A(_01641_),
    .B(_01642_),
    .C(_01643_),
    .X(_01645_));
 sky130_fd_sc_hd__and4bb_1 _07578_ (.A_N(_01644_),
    .B_N(_01645_),
    .C(net761),
    .D(net1801),
    .X(_01646_));
 sky130_fd_sc_hd__nand3_1 _07579_ (.A(_01621_),
    .B(_01640_),
    .C(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__a21o_1 _07580_ (.A1(_01621_),
    .A2(_01640_),
    .B1(_01646_),
    .X(_01648_));
 sky130_fd_sc_hd__a21bo_1 _07581_ (.A1(_01641_),
    .A2(_01643_),
    .B1_N(_01642_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_1 _07582_ (.A(net1883),
    .B(net815),
    .Y(_01650_));
 sky130_fd_sc_hd__and3_1 _07583_ (.A(net1883),
    .B(net815),
    .C(_01649_),
    .X(_01651_));
 sky130_fd_sc_hd__xnor2_1 _07584_ (.A(_01649_),
    .B(_01650_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(net2082),
    .B(net1786),
    .Y(_01653_));
 sky130_fd_sc_hd__and3_1 _07586_ (.A(net2082),
    .B(net1786),
    .C(_01652_),
    .X(_01654_));
 sky130_fd_sc_hd__xnor2_1 _07587_ (.A(_01652_),
    .B(_01653_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand3_1 _07588_ (.A(_01647_),
    .B(_01648_),
    .C(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(_01647_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand3_2 _07590_ (.A(_01632_),
    .B(_01639_),
    .C(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__a21o_1 _07591_ (.A1(_01632_),
    .A2(_01639_),
    .B1(_01657_),
    .X(_01659_));
 sky130_fd_sc_hd__o211ai_2 _07592_ (.A1(_01651_),
    .A2(_01654_),
    .B1(_01658_),
    .C1(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_01658_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand3_2 _07594_ (.A(_01635_),
    .B(_01638_),
    .C(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__a21o_1 _07595_ (.A1(_01635_),
    .A2(_01638_),
    .B1(_01661_),
    .X(_01663_));
 sky130_fd_sc_hd__a211o_1 _07596_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_01651_),
    .C1(_01654_),
    .X(_01664_));
 sky130_fd_sc_hd__o2bb2a_1 _07597_ (.A1_N(net761),
    .A2_N(net1801),
    .B1(_01644_),
    .B2(_01645_),
    .X(_01665_));
 sky130_fd_sc_hd__nor2_1 _07598_ (.A(_01646_),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__and4_1 _07599_ (.A(net2082),
    .B(net761),
    .C(net2824),
    .D(net2819),
    .X(_01667_));
 sky130_fd_sc_hd__nand2_1 _07600_ (.A(net740),
    .B(net1737),
    .Y(_01668_));
 sky130_fd_sc_hd__a22o_1 _07601_ (.A1(net1584),
    .A2(net1168),
    .B1(net1118),
    .B2(net2082),
    .X(_01669_));
 sky130_fd_sc_hd__and2b_1 _07602_ (.A_N(_01667_),
    .B(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__a31o_1 _07603_ (.A1(net740),
    .A2(net1737),
    .A3(_01669_),
    .B1(_01667_),
    .X(_01671_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(net2082),
    .B(net815),
    .Y(_01672_));
 sky130_fd_sc_hd__and3_1 _07605_ (.A(net2082),
    .B(net2773),
    .C(_01671_),
    .X(_01673_));
 sky130_fd_sc_hd__xnor2_1 _07606_ (.A(_01671_),
    .B(_01672_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _07607_ (.A(net1974),
    .B(net1786),
    .Y(_01675_));
 sky130_fd_sc_hd__xnor2_1 _07608_ (.A(_01674_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__and2_1 _07609_ (.A(_01666_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__a21o_1 _07610_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_01655_),
    .X(_01678_));
 sky130_fd_sc_hd__nand3_1 _07611_ (.A(_01656_),
    .B(_01677_),
    .C(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__a31o_1 _07612_ (.A1(net1974),
    .A2(net1786),
    .A3(_01674_),
    .B1(_01673_),
    .X(_01680_));
 sky130_fd_sc_hd__a21o_1 _07613_ (.A1(_01656_),
    .A2(_01678_),
    .B1(_01677_),
    .X(_01681_));
 sky130_fd_sc_hd__nand3_1 _07614_ (.A(_01679_),
    .B(_01680_),
    .C(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _07615_ (.A(_01679_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__and3_1 _07616_ (.A(_01660_),
    .B(_01664_),
    .C(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__a21oi_1 _07617_ (.A1(_01660_),
    .A2(_01664_),
    .B1(_01683_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21o_1 _07618_ (.A1(_01679_),
    .A2(_01681_),
    .B1(_01680_),
    .X(_01686_));
 sky130_fd_sc_hd__xnor2_1 _07619_ (.A(_01668_),
    .B(_01670_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _07620_ (.A(net1974),
    .B(net815),
    .Y(_01688_));
 sky130_fd_sc_hd__and4_1 _07621_ (.A(net1974),
    .B(net761),
    .C(net1737),
    .D(net1118),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _07622_ (.A0(_01688_),
    .A1(net815),
    .S(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__nand2_1 _07623_ (.A(net1694),
    .B(net1786),
    .Y(_01691_));
 sky130_fd_sc_hd__xor2_1 _07624_ (.A(_01690_),
    .B(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_01687_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__xnor2_1 _07626_ (.A(_01666_),
    .B(_01676_),
    .Y(_01694_));
 sky130_fd_sc_hd__nor2_1 _07627_ (.A(_01693_),
    .B(_01694_),
    .Y(_01695_));
 sky130_fd_sc_hd__o2bb2ai_1 _07628_ (.A1_N(net815),
    .A2_N(_01689_),
    .B1(_01690_),
    .B2(_01691_),
    .Y(_01696_));
 sky130_fd_sc_hd__xor2_1 _07629_ (.A(_01693_),
    .B(_01694_),
    .X(_01697_));
 sky130_fd_sc_hd__a21o_1 _07630_ (.A1(_01696_),
    .A2(_01697_),
    .B1(_01695_),
    .X(_01698_));
 sky130_fd_sc_hd__and3_1 _07631_ (.A(_01682_),
    .B(_01686_),
    .C(_01698_),
    .X(_01699_));
 sky130_fd_sc_hd__nand3_1 _07632_ (.A(_01682_),
    .B(_01686_),
    .C(_01698_),
    .Y(_01700_));
 sky130_fd_sc_hd__a21oi_1 _07633_ (.A1(_01682_),
    .A2(_01686_),
    .B1(_01698_),
    .Y(_01701_));
 sky130_fd_sc_hd__xnor2_1 _07634_ (.A(_01696_),
    .B(_01697_),
    .Y(_01702_));
 sky130_fd_sc_hd__or2_1 _07635_ (.A(_01687_),
    .B(_01692_),
    .X(_01703_));
 sky130_fd_sc_hd__and2_1 _07636_ (.A(_01693_),
    .B(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__and4_1 _07637_ (.A(net1694),
    .B(net740),
    .C(net1786),
    .D(net815),
    .X(_01705_));
 sky130_fd_sc_hd__a22oi_1 _07638_ (.A1(net761),
    .A2(net1737),
    .B1(net1118),
    .B2(net1974),
    .Y(_01706_));
 sky130_fd_sc_hd__nor2_1 _07639_ (.A(_01689_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__a22o_1 _07640_ (.A1(net740),
    .A2(net1786),
    .B1(net815),
    .B2(net1694),
    .X(_01708_));
 sky130_fd_sc_hd__and2b_1 _07641_ (.A_N(_01705_),
    .B(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__a21o_1 _07642_ (.A1(_01707_),
    .A2(_01708_),
    .B1(_01705_),
    .X(_01710_));
 sky130_fd_sc_hd__xnor2_1 _07643_ (.A(_01704_),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__xnor2_1 _07644_ (.A(_01707_),
    .B(_01709_),
    .Y(_01712_));
 sky130_fd_sc_hd__and4_1 _07645_ (.A(net740),
    .B(net761),
    .C(net1786),
    .D(net815),
    .X(_01713_));
 sky130_fd_sc_hd__nand2_1 _07646_ (.A(net1694),
    .B(net1118),
    .Y(_01714_));
 sky130_fd_sc_hd__a22o_1 _07647_ (.A1(net761),
    .A2(net1786),
    .B1(net815),
    .B2(net740),
    .X(_01715_));
 sky130_fd_sc_hd__and2b_1 _07648_ (.A_N(_01713_),
    .B(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__a31o_1 _07649_ (.A1(net1694),
    .A2(net1118),
    .A3(_01715_),
    .B1(_01713_),
    .X(_01717_));
 sky130_fd_sc_hd__nand2b_1 _07650_ (.A_N(_01712_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xnor2_1 _07651_ (.A(_01714_),
    .B(_01716_),
    .Y(_01719_));
 sky130_fd_sc_hd__and4_1 _07652_ (.A(net740),
    .B(net761),
    .C(net815),
    .D(net1118),
    .X(_01720_));
 sky130_fd_sc_hd__and2_1 _07653_ (.A(_01719_),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__inv_2 _07654_ (.A(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2b_1 _07655_ (.A_N(_01717_),
    .B(_01712_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(_01718_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__or2_1 _07657_ (.A(_01722_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__a21o_1 _07658_ (.A1(_01718_),
    .A2(_01725_),
    .B1(_01711_),
    .X(_01726_));
 sky130_fd_sc_hd__a21boi_1 _07659_ (.A1(_01704_),
    .A2(_01710_),
    .B1_N(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__nor2_1 _07660_ (.A(_01702_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__or4_2 _07661_ (.A(_01699_),
    .B(_01701_),
    .C(_01702_),
    .D(_01727_),
    .X(_01729_));
 sky130_fd_sc_hd__a211oi_2 _07662_ (.A1(net2777),
    .A2(_01729_),
    .B1(_01684_),
    .C1(_01685_),
    .Y(_01730_));
 sky130_fd_sc_hd__o211ai_2 _07663_ (.A1(_01684_),
    .A2(_01730_),
    .B1(_01662_),
    .C1(_01663_),
    .Y(_01731_));
 sky130_fd_sc_hd__a211oi_1 _07664_ (.A1(_01662_),
    .A2(_01731_),
    .B1(_01636_),
    .C1(_01637_),
    .Y(_01732_));
 sky130_fd_sc_hd__o21ai_1 _07665_ (.A1(_01636_),
    .A2(_01732_),
    .B1(_01610_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _07666_ (.A1(_01609_),
    .A2(_01733_),
    .B1(_01577_),
    .Y(_01734_));
 sky130_fd_sc_hd__o21a_1 _07667_ (.A1(_01575_),
    .A2(_01734_),
    .B1(_01548_),
    .X(_01735_));
 sky130_fd_sc_hd__nor2_1 _07668_ (.A(_01546_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__o21ai_1 _07669_ (.A1(_01546_),
    .A2(_01735_),
    .B1(_01522_),
    .Y(_01737_));
 sky130_fd_sc_hd__xor2_2 _07670_ (.A(_01522_),
    .B(_01736_),
    .X(_01738_));
 sky130_fd_sc_hd__and2b_1 _07671_ (.A_N(_01738_),
    .B(_01464_),
    .X(_01739_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(net1492),
    .B(net1817),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(net1541),
    .B(net758),
    .Y(_01741_));
 sky130_fd_sc_hd__and4_2 _07674_ (.A(net1541),
    .B(net950),
    .C(net1147),
    .D(net758),
    .X(_01742_));
 sky130_fd_sc_hd__nand4_4 _07675_ (.A(net950),
    .B(net818),
    .C(net1147),
    .D(net758),
    .Y(_01743_));
 sky130_fd_sc_hd__a22o_1 _07676_ (.A1(net950),
    .A2(net1147),
    .B1(net758),
    .B2(net1541),
    .X(_01744_));
 sky130_fd_sc_hd__xor2_1 _07677_ (.A(_01742_),
    .B(_01743_),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _07678_ (.A(_01744_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__xor2_1 _07679_ (.A(_01740_),
    .B(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__and4_1 _07680_ (.A(net818),
    .B(net2311),
    .C(net1147),
    .D(net758),
    .X(_01748_));
 sky130_fd_sc_hd__and2_1 _07681_ (.A(_01743_),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__nand2_1 _07682_ (.A(net1541),
    .B(net1817),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _07683_ (.A(_01743_),
    .B(_01748_),
    .Y(_01751_));
 sky130_fd_sc_hd__a22oi_2 _07684_ (.A1(net818),
    .A2(net1147),
    .B1(net758),
    .B2(net950),
    .Y(_01752_));
 sky130_fd_sc_hd__nor4_1 _07685_ (.A(_01749_),
    .B(_01750_),
    .C(_01751_),
    .D(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__o21ai_1 _07686_ (.A1(_01749_),
    .A2(_01753_),
    .B1(_01747_),
    .Y(_01754_));
 sky130_fd_sc_hd__or3_1 _07687_ (.A(_01747_),
    .B(_01749_),
    .C(_01753_),
    .X(_01755_));
 sky130_fd_sc_hd__and2_1 _07688_ (.A(_01754_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__o31a_1 _07689_ (.A1(_01749_),
    .A2(_01751_),
    .A3(_01752_),
    .B1(_01750_),
    .X(_01757_));
 sky130_fd_sc_hd__nor2_1 _07690_ (.A(_01753_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand4_2 _07691_ (.A(net2311),
    .B(net989),
    .C(net1147),
    .D(net758),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_1 _07692_ (.A(_01748_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__nand2_1 _07693_ (.A(net950),
    .B(net1817),
    .Y(_01761_));
 sky130_fd_sc_hd__and2_1 _07694_ (.A(_01748_),
    .B(_01759_),
    .X(_01762_));
 sky130_fd_sc_hd__a22o_1 _07695_ (.A1(net2311),
    .A2(net1147),
    .B1(net758),
    .B2(net818),
    .X(_01763_));
 sky130_fd_sc_hd__or3b_1 _07696_ (.A(_01760_),
    .B(_01762_),
    .C_N(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__nor2_1 _07697_ (.A(_01761_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__o21a_1 _07698_ (.A1(_01760_),
    .A2(_01765_),
    .B1(_01758_),
    .X(_01766_));
 sky130_fd_sc_hd__nor3_1 _07699_ (.A(_01758_),
    .B(_01760_),
    .C(_01765_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _07700_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__and3_1 _07701_ (.A(net1492),
    .B(net1849),
    .C(_01768_),
    .X(_01769_));
 sky130_fd_sc_hd__o21ai_1 _07702_ (.A1(_01766_),
    .A2(_01769_),
    .B1(_01756_),
    .Y(_01770_));
 sky130_fd_sc_hd__or3_1 _07703_ (.A(_01756_),
    .B(_01766_),
    .C(_01769_),
    .X(_01771_));
 sky130_fd_sc_hd__and2_1 _07704_ (.A(_01770_),
    .B(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__a21oi_1 _07705_ (.A1(net1492),
    .A2(net1849),
    .B1(_01768_),
    .Y(_01773_));
 sky130_fd_sc_hd__or2_1 _07706_ (.A(_01769_),
    .B(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__xor2_1 _07707_ (.A(_01761_),
    .B(_01764_),
    .X(_01775_));
 sky130_fd_sc_hd__and4_1 _07708_ (.A(net989),
    .B(net1946),
    .C(net1147),
    .D(net758),
    .X(_01776_));
 sky130_fd_sc_hd__and2_1 _07709_ (.A(_01759_),
    .B(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__a22oi_1 _07710_ (.A1(net818),
    .A2(net1817),
    .B1(net908),
    .B2(net1492),
    .Y(_01778_));
 sky130_fd_sc_hd__and4_1 _07711_ (.A(net1492),
    .B(net818),
    .C(net1817),
    .D(net908),
    .X(_01779_));
 sky130_fd_sc_hd__or2_1 _07712_ (.A(_01778_),
    .B(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__nor2_1 _07713_ (.A(_01759_),
    .B(_01776_),
    .Y(_01781_));
 sky130_fd_sc_hd__a22o_1 _07714_ (.A1(net989),
    .A2(net1147),
    .B1(net758),
    .B2(net2311),
    .X(_01782_));
 sky130_fd_sc_hd__or3b_1 _07715_ (.A(_01777_),
    .B(_01781_),
    .C_N(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__nor2_1 _07716_ (.A(_01780_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o21ai_1 _07717_ (.A1(_01777_),
    .A2(_01784_),
    .B1(_01775_),
    .Y(_01785_));
 sky130_fd_sc_hd__or3_1 _07718_ (.A(_01775_),
    .B(_01777_),
    .C(_01784_),
    .X(_01786_));
 sky130_fd_sc_hd__and2_1 _07719_ (.A(_01785_),
    .B(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__and2_1 _07720_ (.A(net1541),
    .B(net1849),
    .X(_01788_));
 sky130_fd_sc_hd__nor2_1 _07721_ (.A(_01779_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__and2_1 _07722_ (.A(_01779_),
    .B(_01788_),
    .X(_01790_));
 sky130_fd_sc_hd__nor2_1 _07723_ (.A(_01789_),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _07724_ (.A(net1492),
    .B(net2307),
    .Y(_01792_));
 sky130_fd_sc_hd__xnor2_1 _07725_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _07726_ (.A(_01787_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21oi_1 _07727_ (.A1(_01785_),
    .A2(_01794_),
    .B1(_01774_),
    .Y(_01795_));
 sky130_fd_sc_hd__and3_1 _07728_ (.A(_01774_),
    .B(_01785_),
    .C(_01794_),
    .X(_01796_));
 sky130_fd_sc_hd__or2_1 _07729_ (.A(_01795_),
    .B(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__a31o_1 _07730_ (.A1(net1492),
    .A2(net2307),
    .A3(_01791_),
    .B1(_01790_),
    .X(_01798_));
 sky130_fd_sc_hd__and2b_1 _07731_ (.A_N(_01797_),
    .B(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__o21ai_1 _07732_ (.A1(_01795_),
    .A2(_01799_),
    .B1(_01772_),
    .Y(_01800_));
 sky130_fd_sc_hd__or3_1 _07733_ (.A(_01772_),
    .B(_01795_),
    .C(_01799_),
    .X(_01801_));
 sky130_fd_sc_hd__and2_1 _07734_ (.A(_01800_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__and2b_1 _07735_ (.A_N(_01798_),
    .B(_01797_),
    .X(_01803_));
 sky130_fd_sc_hd__or2_1 _07736_ (.A(_01799_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__or2_1 _07737_ (.A(_01787_),
    .B(_01793_),
    .X(_01805_));
 sky130_fd_sc_hd__nand2_1 _07738_ (.A(_01794_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__xnor2_1 _07739_ (.A(_01780_),
    .B(_01783_),
    .Y(_01807_));
 sky130_fd_sc_hd__a22oi_1 _07740_ (.A1(net1946),
    .A2(net1147),
    .B1(net1705),
    .B2(net1960),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_1 _07741_ (.A(_01776_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand4_1 _07742_ (.A(net1492),
    .B(net1636),
    .C(net1147),
    .D(net139),
    .Y(_01810_));
 sky130_fd_sc_hd__and2_1 _07743_ (.A(net1946),
    .B(net1703),
    .X(_01811_));
 sky130_fd_sc_hd__a22o_1 _07744_ (.A1(net1636),
    .A2(net1147),
    .B1(net139),
    .B2(net1492),
    .X(_01812_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_01810_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21bo_1 _07746_ (.A1(_01811_),
    .A2(_01812_),
    .B1_N(_01810_),
    .X(_01814_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_01809_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__or2_1 _07748_ (.A(_01809_),
    .B(_01814_),
    .X(_01816_));
 sky130_fd_sc_hd__and2_1 _07749_ (.A(_01815_),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__a22oi_1 _07750_ (.A1(net2311),
    .A2(net1817),
    .B1(net749),
    .B2(net1492),
    .Y(_01818_));
 sky130_fd_sc_hd__and4_1 _07751_ (.A(net1492),
    .B(net2311),
    .C(net1817),
    .D(net749),
    .X(_01819_));
 sky130_fd_sc_hd__nor2_1 _07752_ (.A(_01818_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _07753_ (.A(net1541),
    .B(net908),
    .Y(_01821_));
 sky130_fd_sc_hd__xor2_1 _07754_ (.A(_01820_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__inv_2 _07755_ (.A(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _07756_ (.A(_01817_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__a21o_1 _07757_ (.A1(_01815_),
    .A2(_01824_),
    .B1(_01807_),
    .X(_01825_));
 sky130_fd_sc_hd__nand3_1 _07758_ (.A(_01807_),
    .B(_01815_),
    .C(_01824_),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_1 _07759_ (.A(_01825_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a31o_1 _07760_ (.A1(net1541),
    .A2(net908),
    .A3(_01820_),
    .B1(_01819_),
    .X(_01828_));
 sky130_fd_sc_hd__a21oi_1 _07761_ (.A1(net1763),
    .A2(net1849),
    .B1(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__and2_1 _07762_ (.A(net1849),
    .B(_01828_),
    .X(_01830_));
 sky130_fd_sc_hd__a21oi_1 _07763_ (.A1(net1761),
    .A2(_01830_),
    .B1(_01829_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand2_1 _07764_ (.A(net1541),
    .B(net2307),
    .Y(_01832_));
 sky130_fd_sc_hd__xor2_1 _07765_ (.A(_01831_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__or2_1 _07766_ (.A(_01827_),
    .B(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__a21o_1 _07767_ (.A1(_01825_),
    .A2(_01834_),
    .B1(_01806_),
    .X(_01835_));
 sky130_fd_sc_hd__nand3_1 _07768_ (.A(_01806_),
    .B(_01825_),
    .C(_01834_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_01835_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__a32o_1 _07770_ (.A1(net1541),
    .A2(net2307),
    .A3(_01831_),
    .B1(_01830_),
    .B2(net1763),
    .X(_01838_));
 sky130_fd_sc_hd__nand2b_1 _07771_ (.A_N(_01837_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21oi_1 _07772_ (.A1(_01835_),
    .A2(_01839_),
    .B1(_01804_),
    .Y(_01840_));
 sky130_fd_sc_hd__and3_1 _07773_ (.A(_01804_),
    .B(_01835_),
    .C(_01839_),
    .X(_01841_));
 sky130_fd_sc_hd__or2_1 _07774_ (.A(_01840_),
    .B(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__xor2_1 _07775_ (.A(_01837_),
    .B(_01838_),
    .X(_01843_));
 sky130_fd_sc_hd__xor2_1 _07776_ (.A(_01827_),
    .B(_01833_),
    .X(_01844_));
 sky130_fd_sc_hd__xnor2_1 _07777_ (.A(_01817_),
    .B(_01823_),
    .Y(_01845_));
 sky130_fd_sc_hd__xnor2_1 _07778_ (.A(_01811_),
    .B(_01813_),
    .Y(_01846_));
 sky130_fd_sc_hd__and4_1 _07779_ (.A(net1541),
    .B(net1636),
    .C(net1705),
    .D(net139),
    .X(_01847_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(_01846_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__xnor2_1 _07781_ (.A(_01846_),
    .B(_01847_),
    .Y(_01849_));
 sky130_fd_sc_hd__a22oi_1 _07782_ (.A1(net1960),
    .A2(net1817),
    .B1(net749),
    .B2(net1541),
    .Y(_01850_));
 sky130_fd_sc_hd__and4_1 _07783_ (.A(net1541),
    .B(net1960),
    .C(net1817),
    .D(net749),
    .X(_01851_));
 sky130_fd_sc_hd__nor2_1 _07784_ (.A(_01850_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(net1763),
    .B(net908),
    .Y(_01853_));
 sky130_fd_sc_hd__xor2_1 _07786_ (.A(_01852_),
    .B(_01853_),
    .X(_01854_));
 sky130_fd_sc_hd__or2_1 _07787_ (.A(_01849_),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__a21oi_1 _07788_ (.A1(_01848_),
    .A2(_01855_),
    .B1(_01845_),
    .Y(_01856_));
 sky130_fd_sc_hd__and3_1 _07789_ (.A(_01845_),
    .B(_01848_),
    .C(_01855_),
    .X(_01857_));
 sky130_fd_sc_hd__or2_1 _07790_ (.A(_01856_),
    .B(_01857_),
    .X(_01858_));
 sky130_fd_sc_hd__a31o_1 _07791_ (.A1(net1763),
    .A2(net908),
    .A3(_01852_),
    .B1(_01851_),
    .X(_01859_));
 sky130_fd_sc_hd__a21oi_1 _07792_ (.A1(net1664),
    .A2(net1849),
    .B1(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__and3_1 _07793_ (.A(net1662),
    .B(net1849),
    .C(_01859_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _07794_ (.A(_01860_),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__a21oi_1 _07795_ (.A1(net1763),
    .A2(net2307),
    .B1(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__and3_1 _07796_ (.A(net1763),
    .B(net2307),
    .C(_01862_),
    .X(_01864_));
 sky130_fd_sc_hd__nor2_1 _07797_ (.A(_01863_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__and2b_1 _07798_ (.A_N(_01858_),
    .B(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__o21ai_1 _07799_ (.A1(_01856_),
    .A2(_01866_),
    .B1(_01844_),
    .Y(_01867_));
 sky130_fd_sc_hd__or3_1 _07800_ (.A(_01844_),
    .B(_01856_),
    .C(_01866_),
    .X(_01868_));
 sky130_fd_sc_hd__and2_1 _07801_ (.A(_01867_),
    .B(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__or2_1 _07802_ (.A(_01861_),
    .B(_01864_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_01869_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21o_1 _07804_ (.A1(_01867_),
    .A2(_01871_),
    .B1(_01843_),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_1 _07805_ (.A(_01843_),
    .B(_01867_),
    .C(_01871_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(_01872_),
    .B(net3459),
    .Y(_01874_));
 sky130_fd_sc_hd__xnor2_1 _07807_ (.A(_01869_),
    .B(_01870_),
    .Y(_01875_));
 sky130_fd_sc_hd__xnor2_1 _07808_ (.A(_01858_),
    .B(_01865_),
    .Y(_01876_));
 sky130_fd_sc_hd__xor2_1 _07809_ (.A(_01849_),
    .B(_01854_),
    .X(_01877_));
 sky130_fd_sc_hd__a22oi_1 _07810_ (.A1(net1636),
    .A2(net1705),
    .B1(net139),
    .B2(net1541),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(_01847_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(net1664),
    .B(net908),
    .Y(_01880_));
 sky130_fd_sc_hd__a22oi_1 _07813_ (.A1(net1946),
    .A2(net1817),
    .B1(net749),
    .B2(net1763),
    .Y(_01881_));
 sky130_fd_sc_hd__and4_1 _07814_ (.A(net1763),
    .B(net1946),
    .C(net1817),
    .D(net749),
    .X(_01882_));
 sky130_fd_sc_hd__nor2_1 _07815_ (.A(_01881_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__xnor2_1 _07816_ (.A(_01880_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__and2_1 _07817_ (.A(_01879_),
    .B(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__nand2_1 _07818_ (.A(_01877_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__xnor2_1 _07819_ (.A(_01877_),
    .B(_01885_),
    .Y(_01887_));
 sky130_fd_sc_hd__a31o_1 _07820_ (.A1(net1664),
    .A2(net908),
    .A3(_01883_),
    .B1(_01882_),
    .X(_01888_));
 sky130_fd_sc_hd__and2_1 _07821_ (.A(net2311),
    .B(net1849),
    .X(_01889_));
 sky130_fd_sc_hd__nor2_1 _07822_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__and2_1 _07823_ (.A(_01888_),
    .B(_01889_),
    .X(_01891_));
 sky130_fd_sc_hd__nor2_1 _07824_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__nand2_1 _07825_ (.A(net1664),
    .B(net2307),
    .Y(_01893_));
 sky130_fd_sc_hd__xor2_1 _07826_ (.A(_01892_),
    .B(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__o21a_1 _07827_ (.A1(_01887_),
    .A2(_01894_),
    .B1(_01886_),
    .X(_01895_));
 sky130_fd_sc_hd__nand2b_1 _07828_ (.A_N(_01895_),
    .B(_01876_),
    .Y(_01896_));
 sky130_fd_sc_hd__xnor2_1 _07829_ (.A(_01876_),
    .B(_01895_),
    .Y(_01897_));
 sky130_fd_sc_hd__o21ba_1 _07830_ (.A1(_01890_),
    .A2(_01893_),
    .B1_N(_01891_),
    .X(_01898_));
 sky130_fd_sc_hd__nand2b_1 _07831_ (.A_N(_01898_),
    .B(_01897_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(_01896_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2b_1 _07833_ (.A_N(_01875_),
    .B(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__xor2_1 _07834_ (.A(_01875_),
    .B(_01900_),
    .X(_01902_));
 sky130_fd_sc_hd__xnor2_1 _07835_ (.A(_01897_),
    .B(_01898_),
    .Y(_01903_));
 sky130_fd_sc_hd__xor2_1 _07836_ (.A(_01887_),
    .B(_01894_),
    .X(_01904_));
 sky130_fd_sc_hd__xnor2_1 _07837_ (.A(_01879_),
    .B(_01884_),
    .Y(_01905_));
 sky130_fd_sc_hd__a22o_1 _07838_ (.A1(net1636),
    .A2(net1817),
    .B1(net749),
    .B2(net1664),
    .X(_01906_));
 sky130_fd_sc_hd__nand4_2 _07839_ (.A(net1664),
    .B(net1636),
    .C(net1817),
    .D(net749),
    .Y(_01907_));
 sky130_fd_sc_hd__and2_1 _07840_ (.A(net2311),
    .B(net908),
    .X(_01908_));
 sky130_fd_sc_hd__a21o_1 _07841_ (.A1(_01906_),
    .A2(_01907_),
    .B1(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__nand3_1 _07842_ (.A(_01906_),
    .B(_01907_),
    .C(_01908_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand4_2 _07843_ (.A(net1763),
    .B(net139),
    .C(_01909_),
    .D(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _07844_ (.A(_01905_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__xor2_1 _07845_ (.A(_01905_),
    .B(_01911_),
    .X(_01913_));
 sky130_fd_sc_hd__a21bo_1 _07846_ (.A1(_01906_),
    .A2(_01908_),
    .B1_N(_01907_),
    .X(_01914_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(net1960),
    .B(net1849),
    .Y(_01915_));
 sky130_fd_sc_hd__and3_1 _07848_ (.A(net1960),
    .B(net1849),
    .C(_01914_),
    .X(_01916_));
 sky130_fd_sc_hd__xnor2_1 _07849_ (.A(_01914_),
    .B(_01915_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _07850_ (.A(net2311),
    .B(net2307),
    .Y(_01918_));
 sky130_fd_sc_hd__xor2_1 _07851_ (.A(_01917_),
    .B(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__inv_2 _07852_ (.A(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__a21oi_1 _07853_ (.A1(_01913_),
    .A2(_01920_),
    .B1(_01912_),
    .Y(_01921_));
 sky130_fd_sc_hd__and2b_1 _07854_ (.A_N(_01921_),
    .B(_01904_),
    .X(_01922_));
 sky130_fd_sc_hd__xnor2_1 _07855_ (.A(_01904_),
    .B(_01921_),
    .Y(_01923_));
 sky130_fd_sc_hd__a31oi_2 _07856_ (.A1(net2311),
    .A2(net2307),
    .A3(_01917_),
    .B1(_01916_),
    .Y(_01924_));
 sky130_fd_sc_hd__and2b_1 _07857_ (.A_N(_01924_),
    .B(_01923_),
    .X(_01925_));
 sky130_fd_sc_hd__nor2_1 _07858_ (.A(_01922_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2b_1 _07859_ (.A_N(_01926_),
    .B(_01903_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_1 _07860_ (.A(_01903_),
    .B(_01926_),
    .Y(_01928_));
 sky130_fd_sc_hd__xnor2_1 _07861_ (.A(_01923_),
    .B(_01924_),
    .Y(_01929_));
 sky130_fd_sc_hd__xnor2_1 _07862_ (.A(_01913_),
    .B(_01920_),
    .Y(_01930_));
 sky130_fd_sc_hd__a22o_1 _07863_ (.A1(net1763),
    .A2(net139),
    .B1(_01909_),
    .B2(_01910_),
    .X(_01931_));
 sky130_fd_sc_hd__a22o_1 _07864_ (.A1(net1960),
    .A2(net908),
    .B1(net749),
    .B2(net2311),
    .X(_01932_));
 sky130_fd_sc_hd__and4_1 _07865_ (.A(net2311),
    .B(net1960),
    .C(net908),
    .D(net749),
    .X(_01933_));
 sky130_fd_sc_hd__nand4_1 _07866_ (.A(net2311),
    .B(net1960),
    .C(net908),
    .D(net749),
    .Y(_01934_));
 sky130_fd_sc_hd__and4_1 _07867_ (.A(net1664),
    .B(net139),
    .C(_01932_),
    .D(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nand4_1 _07868_ (.A(net1664),
    .B(net139),
    .C(_01932_),
    .D(_01934_),
    .Y(_01936_));
 sky130_fd_sc_hd__nand3_1 _07869_ (.A(_01911_),
    .B(_01931_),
    .C(_01935_),
    .Y(_01937_));
 sky130_fd_sc_hd__a21o_1 _07870_ (.A1(_01911_),
    .A2(_01931_),
    .B1(_01935_),
    .X(_01938_));
 sky130_fd_sc_hd__a21oi_1 _07871_ (.A1(net1946),
    .A2(net1849),
    .B1(_01933_),
    .Y(_01939_));
 sky130_fd_sc_hd__and3_1 _07872_ (.A(net1946),
    .B(net1849),
    .C(_01933_),
    .X(_01940_));
 sky130_fd_sc_hd__or2_1 _07873_ (.A(_01939_),
    .B(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_1 _07874_ (.A(net1960),
    .B(net2307),
    .Y(_01942_));
 sky130_fd_sc_hd__xor2_1 _07875_ (.A(_01941_),
    .B(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__nand3_1 _07876_ (.A(_01937_),
    .B(_01938_),
    .C(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__and2_1 _07877_ (.A(_01937_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__nor2_1 _07878_ (.A(_01930_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__xnor2_1 _07879_ (.A(_01930_),
    .B(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__o21ba_1 _07880_ (.A1(_01939_),
    .A2(_01942_),
    .B1_N(_01940_),
    .X(_01948_));
 sky130_fd_sc_hd__o21ba_1 _07881_ (.A1(_01947_),
    .A2(_01948_),
    .B1_N(_01946_),
    .X(_01949_));
 sky130_fd_sc_hd__and2b_1 _07882_ (.A_N(_01949_),
    .B(_01929_),
    .X(_01950_));
 sky130_fd_sc_hd__xnor2_1 _07883_ (.A(_01929_),
    .B(_01949_),
    .Y(_01951_));
 sky130_fd_sc_hd__xnor2_1 _07884_ (.A(_01947_),
    .B(_01948_),
    .Y(_01952_));
 sky130_fd_sc_hd__a21o_1 _07885_ (.A1(_01937_),
    .A2(_01938_),
    .B1(_01943_),
    .X(_01953_));
 sky130_fd_sc_hd__a22o_1 _07886_ (.A1(net1664),
    .A2(net139),
    .B1(_01932_),
    .B2(_01934_),
    .X(_01954_));
 sky130_fd_sc_hd__a22o_1 _07887_ (.A1(net1946),
    .A2(net908),
    .B1(net749),
    .B2(net1960),
    .X(_01955_));
 sky130_fd_sc_hd__nand4_2 _07888_ (.A(net1958),
    .B(net1946),
    .C(net2499),
    .D(net749),
    .Y(_01956_));
 sky130_fd_sc_hd__and4_1 _07889_ (.A(net2311),
    .B(net139),
    .C(_01955_),
    .D(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__and3_1 _07890_ (.A(_01936_),
    .B(_01954_),
    .C(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__a21o_1 _07891_ (.A1(_01936_),
    .A2(_01954_),
    .B1(_01957_),
    .X(_01959_));
 sky130_fd_sc_hd__nand2b_1 _07892_ (.A_N(_01958_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__nand2_1 _07893_ (.A(net1636),
    .B(net1849),
    .Y(_01961_));
 sky130_fd_sc_hd__xnor2_1 _07894_ (.A(_01956_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(net1946),
    .B(net2307),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _07896_ (.A(_01962_),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _07897_ (.A(_01962_),
    .B(_01963_),
    .X(_01965_));
 sky130_fd_sc_hd__and2_1 _07898_ (.A(_01964_),
    .B(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__a21o_1 _07899_ (.A1(_01959_),
    .A2(_01966_),
    .B1(_01958_),
    .X(_01967_));
 sky130_fd_sc_hd__nand3_1 _07900_ (.A(_01944_),
    .B(_01953_),
    .C(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__a21o_1 _07901_ (.A1(_01944_),
    .A2(_01953_),
    .B1(_01967_),
    .X(_01969_));
 sky130_fd_sc_hd__o21ai_1 _07902_ (.A1(_01956_),
    .A2(_01961_),
    .B1(_01965_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand3_1 _07903_ (.A(_01968_),
    .B(_01969_),
    .C(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _07904_ (.A(_01968_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__and2b_1 _07905_ (.A_N(_01952_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__a21o_1 _07906_ (.A1(_01968_),
    .A2(_01969_),
    .B1(_01970_),
    .X(_01974_));
 sky130_fd_sc_hd__xnor2_2 _07907_ (.A(_01960_),
    .B(_01966_),
    .Y(_01975_));
 sky130_fd_sc_hd__a22oi_1 _07908_ (.A1(net2311),
    .A2(net139),
    .B1(_01955_),
    .B2(_01956_),
    .Y(_01976_));
 sky130_fd_sc_hd__or2_1 _07909_ (.A(_01957_),
    .B(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_1 _07910_ (.A1(net1636),
    .A2(net2499),
    .B1(net749),
    .B2(net1946),
    .X(_01978_));
 sky130_fd_sc_hd__and3_1 _07911_ (.A(net1946),
    .B(net1636),
    .C(net2534),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _07912_ (.A(net908),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__nand4_2 _07913_ (.A(net1960),
    .B(net1361),
    .C(_01978_),
    .D(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__or2_1 _07914_ (.A(_01977_),
    .B(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__xnor2_2 _07915_ (.A(_01977_),
    .B(_01981_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _07916_ (.A(net1636),
    .B(net2307),
    .Y(_01984_));
 sky130_fd_sc_hd__nand3_1 _07917_ (.A(net2307),
    .B(net908),
    .C(_01979_),
    .Y(_01985_));
 sky130_fd_sc_hd__a21bo_1 _07918_ (.A1(_01980_),
    .A2(_01984_),
    .B1_N(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__o21ai_2 _07919_ (.A1(_01983_),
    .A2(_01986_),
    .B1(_01982_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand2_1 _07920_ (.A(_01975_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _07921_ (.A(_01975_),
    .B(_01987_),
    .Y(_01989_));
 sky130_fd_sc_hd__xor2_1 _07922_ (.A(_01975_),
    .B(_01987_),
    .X(_01990_));
 sky130_fd_sc_hd__o21ai_1 _07923_ (.A1(_01985_),
    .A2(_01989_),
    .B1(_01988_),
    .Y(_01991_));
 sky130_fd_sc_hd__and3_1 _07924_ (.A(_01971_),
    .B(_01974_),
    .C(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__a21oi_1 _07925_ (.A1(_01971_),
    .A2(_01974_),
    .B1(_01991_),
    .Y(_01993_));
 sky130_fd_sc_hd__xnor2_1 _07926_ (.A(_01985_),
    .B(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__xor2_1 _07927_ (.A(_01983_),
    .B(_01986_),
    .X(_01995_));
 sky130_fd_sc_hd__a22o_1 _07928_ (.A1(net1960),
    .A2(net139),
    .B1(_01978_),
    .B2(_01980_),
    .X(_01996_));
 sky130_fd_sc_hd__and2_1 _07929_ (.A(net139),
    .B(_01979_),
    .X(_01997_));
 sky130_fd_sc_hd__and3_1 _07930_ (.A(_01981_),
    .B(_01996_),
    .C(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__and2_1 _07931_ (.A(_01995_),
    .B(_01998_),
    .X(_01999_));
 sky130_fd_sc_hd__and4bb_2 _07932_ (.A_N(_01992_),
    .B_N(_01993_),
    .C(_01994_),
    .D(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__xor2_1 _07933_ (.A(_01952_),
    .B(_01972_),
    .X(_02001_));
 sky130_fd_sc_hd__o21ba_1 _07934_ (.A1(_01992_),
    .A2(_02000_),
    .B1_N(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__o21a_1 _07935_ (.A1(_01973_),
    .A2(_02002_),
    .B1(_01951_),
    .X(_02003_));
 sky130_fd_sc_hd__o21ai_1 _07936_ (.A1(_01950_),
    .A2(_02003_),
    .B1(_01928_),
    .Y(_02004_));
 sky130_fd_sc_hd__a21o_1 _07937_ (.A1(_01927_),
    .A2(_02004_),
    .B1(_01902_),
    .X(_02005_));
 sky130_fd_sc_hd__a21o_1 _07938_ (.A1(_01901_),
    .A2(_02005_),
    .B1(_01874_),
    .X(_02006_));
 sky130_fd_sc_hd__a21oi_1 _07939_ (.A1(_01872_),
    .A2(_02006_),
    .B1(_01842_),
    .Y(_02007_));
 sky130_fd_sc_hd__o21ai_1 _07940_ (.A1(_01840_),
    .A2(_02007_),
    .B1(_01802_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(_01800_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__o22ai_4 _07942_ (.A1(_01742_),
    .A2(_01743_),
    .B1(_01746_),
    .B2(_01740_),
    .Y(_02010_));
 sky130_fd_sc_hd__a22o_1 _07943_ (.A1(net1541),
    .A2(net1147),
    .B1(net758),
    .B2(net1492),
    .X(_02011_));
 sky130_fd_sc_hd__nand4_1 _07944_ (.A(net1492),
    .B(net1541),
    .C(net1147),
    .D(net758),
    .Y(_02012_));
 sky130_fd_sc_hd__a21oi_1 _07945_ (.A1(_02011_),
    .A2(_02012_),
    .B1(_01742_),
    .Y(_02013_));
 sky130_fd_sc_hd__and2b_1 _07946_ (.A_N(net1492),
    .B(_01742_),
    .X(_02014_));
 sky130_fd_sc_hd__nor2_1 _07947_ (.A(_02013_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__xnor2_2 _07948_ (.A(_02010_),
    .B(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _07949_ (.A(_01754_),
    .B(_01770_),
    .Y(_02017_));
 sky130_fd_sc_hd__xor2_2 _07950_ (.A(_02016_),
    .B(_02017_),
    .X(_02018_));
 sky130_fd_sc_hd__inv_2 _07951_ (.A(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__xnor2_2 _07952_ (.A(_02009_),
    .B(_02018_),
    .Y(_02020_));
 sky130_fd_sc_hd__xnor2_2 _07953_ (.A(_01464_),
    .B(_01738_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21o_1 _07954_ (.A1(_02020_),
    .A2(_02021_),
    .B1(_01739_),
    .X(_02022_));
 sky130_fd_sc_hd__a2bb2o_1 _07955_ (.A1_N(_01770_),
    .A2_N(_02016_),
    .B1(_02019_),
    .B2(_02009_),
    .X(_02023_));
 sky130_fd_sc_hd__nor2_1 _07956_ (.A(_01754_),
    .B(_02016_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21o_1 _07957_ (.A1(_02010_),
    .A2(_02015_),
    .B1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__a31o_1 _07958_ (.A1(net1492),
    .A2(net1147),
    .A3(_01741_),
    .B1(_02014_),
    .X(_02026_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__or2_1 _07960_ (.A(_02025_),
    .B(_02026_),
    .X(_02028_));
 sky130_fd_sc_hd__and2_1 _07961_ (.A(_02027_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _07962_ (.A(_02023_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__or2_1 _07963_ (.A(_02023_),
    .B(_02029_),
    .X(_02031_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_02030_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__a22o_1 _07965_ (.A1(net1550),
    .A2(net848),
    .B1(net770),
    .B2(net1496),
    .X(_02033_));
 sky130_fd_sc_hd__nand4_1 _07966_ (.A(net1496),
    .B(net1550),
    .C(net848),
    .D(net770),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07967_ (.A(_02033_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21o_1 _07968_ (.A1(_00698_),
    .A2(_00700_),
    .B1(_00703_),
    .X(_02036_));
 sky130_fd_sc_hd__xnor2_1 _07969_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__xnor2_1 _07970_ (.A(_00697_),
    .B(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__a21o_1 _07971_ (.A1(_00716_),
    .A2(_00719_),
    .B1(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__nand3_1 _07972_ (.A(_00716_),
    .B(_00719_),
    .C(_02038_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _07973_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__or2_1 _07974_ (.A(_00739_),
    .B(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__nand2_1 _07975_ (.A(_00739_),
    .B(_02041_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_2 _07976_ (.A(_02042_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21oi_2 _07977_ (.A1(_00767_),
    .A2(_00951_),
    .B1(_00765_),
    .Y(_02045_));
 sky130_fd_sc_hd__xnor2_2 _07978_ (.A(_02044_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__a21o_2 _07979_ (.A1(_01022_),
    .A2(_01209_),
    .B1(_01021_),
    .X(_02047_));
 sky130_fd_sc_hd__o21ba_1 _07980_ (.A1(_00955_),
    .A2(_00961_),
    .B1_N(_00963_),
    .X(_02048_));
 sky130_fd_sc_hd__and4_1 _07981_ (.A(net1456),
    .B(net697),
    .C(net752),
    .D(net2152),
    .X(_02049_));
 sky130_fd_sc_hd__a32o_1 _07982_ (.A1(net1456),
    .A2(net2152),
    .A3(_00956_),
    .B1(net697),
    .B2(net752),
    .X(_02050_));
 sky130_fd_sc_hd__a21bo_1 _07983_ (.A1(_00956_),
    .A2(_02049_),
    .B1_N(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__nor2_1 _07984_ (.A(_02048_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__xnor2_1 _07985_ (.A(_02048_),
    .B(_02051_),
    .Y(_02053_));
 sky130_fd_sc_hd__inv_2 _07986_ (.A(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _07987_ (.A(_00975_),
    .B(_00997_),
    .Y(_02055_));
 sky130_fd_sc_hd__xnor2_1 _07988_ (.A(_02053_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__inv_2 _07989_ (.A(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__xnor2_2 _07990_ (.A(_02047_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _07991_ (.A(_02046_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__a22oi_1 _07992_ (.A1(net725),
    .A2(net1853),
    .B1(net779),
    .B2(net1504),
    .Y(_02060_));
 sky130_fd_sc_hd__and4_1 _07993_ (.A(net1504),
    .B(net725),
    .C(net1853),
    .D(net779),
    .X(_02061_));
 sky130_fd_sc_hd__nor2_1 _07994_ (.A(_02060_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__a32o_1 _07995_ (.A1(net1504),
    .A2(net2114),
    .A3(_01212_),
    .B1(_01213_),
    .B2(net920),
    .X(_02063_));
 sky130_fd_sc_hd__nand2_1 _07996_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__or2_1 _07997_ (.A(_02062_),
    .B(_02063_),
    .X(_02065_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(_01222_),
    .B(_01236_),
    .Y(_02067_));
 sky130_fd_sc_hd__xnor2_1 _08000_ (.A(_02066_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2b_1 _08001_ (.A_N(_01255_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__xnor2_1 _08002_ (.A(_01255_),
    .B(_02068_),
    .Y(_02070_));
 sky130_fd_sc_hd__o21ai_2 _08003_ (.A1(_01280_),
    .A2(_01460_),
    .B1(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__or3_1 _08004_ (.A(_01280_),
    .B(_01460_),
    .C(_02070_),
    .X(_02072_));
 sky130_fd_sc_hd__nand2_1 _08005_ (.A(_02071_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__xor2_2 _08006_ (.A(_02046_),
    .B(_02058_),
    .X(_02074_));
 sky130_fd_sc_hd__a31o_2 _08007_ (.A1(_02071_),
    .A2(_02072_),
    .A3(_02074_),
    .B1(_02059_),
    .X(_02075_));
 sky130_fd_sc_hd__and3_1 _08008_ (.A(net1411),
    .B(net1777),
    .C(_01465_),
    .X(_02076_));
 sky130_fd_sc_hd__o21ai_2 _08009_ (.A1(_01475_),
    .A2(_01518_),
    .B1(_01516_),
    .Y(_02077_));
 sky130_fd_sc_hd__xor2_1 _08010_ (.A(_02076_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_1 _08011_ (.A(_01490_),
    .B(_01518_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _08012_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21oi_1 _08013_ (.A1(_01521_),
    .A2(_01737_),
    .B1(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__and3_1 _08014_ (.A(_01521_),
    .B(_01737_),
    .C(_02080_),
    .X(_02082_));
 sky130_fd_sc_hd__or2_2 _08015_ (.A(_02081_),
    .B(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__and2b_1 _08016_ (.A_N(_02083_),
    .B(_02075_),
    .X(_02084_));
 sky130_fd_sc_hd__xnor2_2 _08017_ (.A(_02075_),
    .B(_02083_),
    .Y(_02085_));
 sky130_fd_sc_hd__and2b_1 _08018_ (.A_N(_02032_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__xor2_2 _08019_ (.A(_02032_),
    .B(_02085_),
    .X(_02087_));
 sky130_fd_sc_hd__and3_1 _08020_ (.A(net1504),
    .B(net1853),
    .C(_01211_),
    .X(_02088_));
 sky130_fd_sc_hd__o21ai_1 _08021_ (.A1(_01222_),
    .A2(_02066_),
    .B1(_02064_),
    .Y(_02089_));
 sky130_fd_sc_hd__xor2_1 _08022_ (.A(_02088_),
    .B(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__nor2_1 _08023_ (.A(_01236_),
    .B(_02066_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(_02090_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__xnor2_1 _08025_ (.A(_02090_),
    .B(_02091_),
    .Y(_02093_));
 sky130_fd_sc_hd__a21o_1 _08026_ (.A1(_02069_),
    .A2(_02071_),
    .B1(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__nand3_1 _08027_ (.A(_02069_),
    .B(_02071_),
    .C(_02093_),
    .Y(_02095_));
 sky130_fd_sc_hd__and2_2 _08028_ (.A(_02094_),
    .B(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__inv_2 _08029_ (.A(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__a32o_1 _08030_ (.A1(_02033_),
    .A2(_02034_),
    .A3(_02036_),
    .B1(_02037_),
    .B2(_00697_),
    .X(_02098_));
 sky130_fd_sc_hd__and3b_1 _08031_ (.A_N(_00695_),
    .B(net848),
    .C(net1496),
    .X(_02099_));
 sky130_fd_sc_hd__and2_1 _08032_ (.A(_02098_),
    .B(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__xor2_2 _08033_ (.A(_02098_),
    .B(_02099_),
    .X(_02101_));
 sky130_fd_sc_hd__and2b_1 _08034_ (.A_N(_02039_),
    .B(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__xnor2_2 _08035_ (.A(_02039_),
    .B(_02101_),
    .Y(_02103_));
 sky130_fd_sc_hd__o21ai_2 _08036_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02042_),
    .Y(_02104_));
 sky130_fd_sc_hd__xor2_2 _08037_ (.A(_02103_),
    .B(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__a22oi_4 _08038_ (.A1(_00997_),
    .A2(_02054_),
    .B1(_02057_),
    .B2(_02047_),
    .Y(_02106_));
 sky130_fd_sc_hd__and2_1 _08039_ (.A(_00975_),
    .B(_02054_),
    .X(_02107_));
 sky130_fd_sc_hd__or2_1 _08040_ (.A(_02052_),
    .B(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__a21o_1 _08041_ (.A1(net1456),
    .A2(net752),
    .B1(_00954_),
    .X(_02109_));
 sky130_fd_sc_hd__and2b_1 _08042_ (.A_N(_02049_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__xnor2_2 _08043_ (.A(_02108_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__xor2_2 _08044_ (.A(_02106_),
    .B(_02111_),
    .X(_02112_));
 sky130_fd_sc_hd__nand2_1 _08045_ (.A(_02105_),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__xnor2_2 _08046_ (.A(_02105_),
    .B(_02112_),
    .Y(_02114_));
 sky130_fd_sc_hd__xor2_2 _08047_ (.A(_02096_),
    .B(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__a22oi_1 _08048_ (.A1(net537),
    .A2(net2686),
    .B1(net1164),
    .B2(net1385),
    .Y(_02116_));
 sky130_fd_sc_hd__and4_1 _08049_ (.A(net1385),
    .B(net537),
    .C(net2686),
    .D(net1164),
    .X(_02117_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_1 _08051_ (.A(net537),
    .B(net1164),
    .Y(_02119_));
 sky130_fd_sc_hd__and4_1 _08052_ (.A(net537),
    .B(net1160),
    .C(net2686),
    .D(net1164),
    .X(_02120_));
 sky130_fd_sc_hd__a22o_1 _08053_ (.A1(net1160),
    .A2(net2686),
    .B1(net1164),
    .B2(net537),
    .X(_02121_));
 sky130_fd_sc_hd__and2b_1 _08054_ (.A_N(_02120_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__nand2_1 _08055_ (.A(net1385),
    .B(net2678),
    .Y(_02123_));
 sky130_fd_sc_hd__a31o_1 _08056_ (.A1(net1385),
    .A2(net2678),
    .A3(_02121_),
    .B1(_02120_),
    .X(_02124_));
 sky130_fd_sc_hd__and2_1 _08057_ (.A(_02118_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__xor2_1 _08058_ (.A(_02122_),
    .B(_02123_),
    .X(_02126_));
 sky130_fd_sc_hd__nand4_1 _08059_ (.A(net1160),
    .B(net2247),
    .C(net2686),
    .D(net1164),
    .Y(_02127_));
 sky130_fd_sc_hd__a22o_1 _08060_ (.A1(net2247),
    .A2(net2686),
    .B1(net1164),
    .B2(net1160),
    .X(_02128_));
 sky130_fd_sc_hd__nand2_1 _08061_ (.A(_02127_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _08062_ (.A(net1480),
    .B(net2678),
    .Y(_02130_));
 sky130_fd_sc_hd__o21ai_1 _08063_ (.A1(_02129_),
    .A2(_02130_),
    .B1(_02127_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand2b_1 _08064_ (.A_N(_02126_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _08065_ (.A(_02118_),
    .B(_02124_),
    .Y(_02133_));
 sky130_fd_sc_hd__or2_2 _08066_ (.A(_02125_),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o21bai_2 _08067_ (.A1(_02132_),
    .A2(_02134_),
    .B1_N(_02125_),
    .Y(_02135_));
 sky130_fd_sc_hd__and3_1 _08068_ (.A(net1385),
    .B(net2686),
    .C(_02119_),
    .X(_02136_));
 sky130_fd_sc_hd__xnor2_2 _08069_ (.A(_02135_),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__inv_2 _08070_ (.A(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2b_1 _08071_ (.A_N(_02131_),
    .B(_02126_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_02132_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__xnor2_2 _08073_ (.A(_02129_),
    .B(_02130_),
    .Y(_02141_));
 sky130_fd_sc_hd__inv_2 _08074_ (.A(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand4_1 _08075_ (.A(net2247),
    .B(net977),
    .C(net1091),
    .D(net2803),
    .Y(_02143_));
 sky130_fd_sc_hd__a22o_1 _08076_ (.A1(net977),
    .A2(net1091),
    .B1(net2803),
    .B2(net2247),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(net1160),
    .B(net2678),
    .Y(_02146_));
 sky130_fd_sc_hd__o21ai_1 _08079_ (.A1(_02145_),
    .A2(_02146_),
    .B1(_02143_),
    .Y(_02147_));
 sky130_fd_sc_hd__xnor2_1 _08080_ (.A(_02141_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__and3_1 _08081_ (.A(net1385),
    .B(net734),
    .C(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__a21oi_1 _08082_ (.A1(_02142_),
    .A2(_02147_),
    .B1(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__or2_1 _08083_ (.A(_02140_),
    .B(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__nor2_2 _08084_ (.A(_02134_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__xnor2_2 _08085_ (.A(_02137_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _08086_ (.A(_02140_),
    .B(_02150_),
    .Y(_02154_));
 sky130_fd_sc_hd__and2_1 _08087_ (.A(_02151_),
    .B(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__a21oi_1 _08088_ (.A1(net1385),
    .A2(net734),
    .B1(_02148_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _08089_ (.A(_02149_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_1 _08090_ (.A(_02145_),
    .B(_02146_),
    .Y(_02158_));
 sky130_fd_sc_hd__and4_1 _08091_ (.A(net977),
    .B(net866),
    .C(net1091),
    .D(net1164),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_1 _08092_ (.A1(net866),
    .A2(net1091),
    .B1(net1164),
    .B2(net977),
    .X(_02160_));
 sky130_fd_sc_hd__nand2b_1 _08093_ (.A_N(_02159_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _08094_ (.A(net2247),
    .B(net1085),
    .Y(_02162_));
 sky130_fd_sc_hd__a31o_1 _08095_ (.A1(net2247),
    .A2(net1085),
    .A3(_02160_),
    .B1(_02159_),
    .X(_02163_));
 sky130_fd_sc_hd__and2b_1 _08096_ (.A_N(_02158_),
    .B(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__and2b_1 _08097_ (.A_N(_02163_),
    .B(_02158_),
    .X(_02165_));
 sky130_fd_sc_hd__or2_1 _08098_ (.A(_02164_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__a22oi_1 _08099_ (.A1(net537),
    .A2(net734),
    .B1(net1176),
    .B2(net1385),
    .Y(_02167_));
 sky130_fd_sc_hd__and4_2 _08100_ (.A(net1385),
    .B(net537),
    .C(net3010),
    .D(net1176),
    .X(_02168_));
 sky130_fd_sc_hd__nor2_1 _08101_ (.A(_02167_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__and2b_1 _08102_ (.A_N(_02166_),
    .B(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__o21a_1 _08103_ (.A1(_02164_),
    .A2(_02170_),
    .B1(_02157_),
    .X(_02171_));
 sky130_fd_sc_hd__nor3_1 _08104_ (.A(_02157_),
    .B(_02164_),
    .C(_02170_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_2 _08105_ (.A(_02171_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__a21oi_1 _08106_ (.A1(_02168_),
    .A2(_02173_),
    .B1(_02171_),
    .Y(_02174_));
 sky130_fd_sc_hd__and2b_1 _08107_ (.A_N(_02174_),
    .B(_02155_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2_1 _08108_ (.A(_02132_),
    .B(_02151_),
    .Y(_02176_));
 sky130_fd_sc_hd__xnor2_1 _08109_ (.A(_02134_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_1 _08110_ (.A(_02175_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__or2_1 _08111_ (.A(_02175_),
    .B(_02177_),
    .X(_02179_));
 sky130_fd_sc_hd__nand2_1 _08112_ (.A(_02178_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__and2b_1 _08113_ (.A_N(_02155_),
    .B(_02174_),
    .X(_02181_));
 sky130_fd_sc_hd__or2_1 _08114_ (.A(_02175_),
    .B(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__xnor2_4 _08115_ (.A(_02168_),
    .B(_02173_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_2 _08116_ (.A(_02166_),
    .B(_02169_),
    .Y(_02184_));
 sky130_fd_sc_hd__xnor2_1 _08117_ (.A(_02161_),
    .B(_02162_),
    .Y(_02185_));
 sky130_fd_sc_hd__and4_1 _08118_ (.A(net866),
    .B(net884),
    .C(net1091),
    .D(net1164),
    .X(_02186_));
 sky130_fd_sc_hd__a22o_1 _08119_ (.A1(net884),
    .A2(net1091),
    .B1(net1164),
    .B2(net1790),
    .X(_02187_));
 sky130_fd_sc_hd__nand2b_1 _08120_ (.A_N(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _08121_ (.A(net977),
    .B(net1085),
    .Y(_02189_));
 sky130_fd_sc_hd__a31o_1 _08122_ (.A1(net2256),
    .A2(net1085),
    .A3(_02187_),
    .B1(_02186_),
    .X(_02190_));
 sky130_fd_sc_hd__and2b_1 _08123_ (.A_N(_02185_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__xor2_1 _08124_ (.A(_02185_),
    .B(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__a22o_1 _08125_ (.A1(net1160),
    .A2(net733),
    .B1(net1176),
    .B2(net537),
    .X(_02193_));
 sky130_fd_sc_hd__and4_1 _08126_ (.A(net537),
    .B(net1160),
    .C(net3010),
    .D(net1176),
    .X(_02194_));
 sky130_fd_sc_hd__nand4_1 _08127_ (.A(net537),
    .B(net1160),
    .C(net734),
    .D(net1175),
    .Y(_02195_));
 sky130_fd_sc_hd__a22oi_1 _08128_ (.A1(net1385),
    .A2(net1082),
    .B1(_02193_),
    .B2(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__and4_1 _08129_ (.A(net1385),
    .B(net1082),
    .C(_02193_),
    .D(_02195_),
    .X(_02197_));
 sky130_fd_sc_hd__or2_1 _08130_ (.A(_02196_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__nor2_1 _08131_ (.A(_02192_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__o21ai_4 _08132_ (.A1(_02191_),
    .A2(_02199_),
    .B1(_02184_),
    .Y(_02200_));
 sky130_fd_sc_hd__or3_2 _08133_ (.A(_02184_),
    .B(_02191_),
    .C(_02199_),
    .X(_02201_));
 sky130_fd_sc_hd__o211ai_4 _08134_ (.A1(_02194_),
    .A2(net3812),
    .B1(_02200_),
    .C1(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_2 _08135_ (.A(_02200_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2b_1 _08136_ (.A_N(_02183_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _08137_ (.A(_02182_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__and2_1 _08138_ (.A(_02182_),
    .B(_02204_),
    .X(_02206_));
 sky130_fd_sc_hd__nor2_1 _08139_ (.A(_02205_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__xor2_4 _08140_ (.A(_02183_),
    .B(_02203_),
    .X(_02208_));
 sky130_fd_sc_hd__a211o_1 _08141_ (.A1(_02200_),
    .A2(_02201_),
    .B1(_02194_),
    .C1(net3812),
    .X(_02209_));
 sky130_fd_sc_hd__xor2_1 _08142_ (.A(_02192_),
    .B(_02198_),
    .X(_02210_));
 sky130_fd_sc_hd__xnor2_1 _08143_ (.A(_02188_),
    .B(_02189_),
    .Y(_02211_));
 sky130_fd_sc_hd__nand4_2 _08144_ (.A(net884),
    .B(net1603),
    .C(net2686),
    .D(net1164),
    .Y(_02212_));
 sky130_fd_sc_hd__a22o_1 _08145_ (.A1(net1603),
    .A2(net1091),
    .B1(net1164),
    .B2(net884),
    .X(_02213_));
 sky130_fd_sc_hd__nand4_1 _08146_ (.A(net866),
    .B(net2678),
    .C(_02212_),
    .D(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(_02212_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__and2b_1 _08148_ (.A_N(_02211_),
    .B(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__a22o_1 _08149_ (.A1(net2247),
    .A2(net734),
    .B1(net1175),
    .B2(net1160),
    .X(_02217_));
 sky130_fd_sc_hd__nand4_1 _08150_ (.A(net1160),
    .B(net2247),
    .C(net734),
    .D(net2970),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_02217_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2_1 _08152_ (.A(net537),
    .B(net1082),
    .Y(_02220_));
 sky130_fd_sc_hd__xnor2_1 _08153_ (.A(_02219_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__xor2_1 _08154_ (.A(_02211_),
    .B(_02215_),
    .X(_02222_));
 sky130_fd_sc_hd__nor2_1 _08155_ (.A(_02221_),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__o21a_1 _08156_ (.A1(_02216_),
    .A2(_02223_),
    .B1(_02210_),
    .X(_02224_));
 sky130_fd_sc_hd__o21ai_1 _08157_ (.A1(_02219_),
    .A2(_02220_),
    .B1(_02218_),
    .Y(_02225_));
 sky130_fd_sc_hd__or3_1 _08158_ (.A(_02210_),
    .B(_02216_),
    .C(_02223_),
    .X(_02226_));
 sky130_fd_sc_hd__nand2b_1 _08159_ (.A_N(_02224_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__and2b_1 _08160_ (.A_N(_02227_),
    .B(_02225_),
    .X(_02228_));
 sky130_fd_sc_hd__o211ai_2 _08161_ (.A1(_02224_),
    .A2(_02228_),
    .B1(_02202_),
    .C1(_02209_),
    .Y(_02229_));
 sky130_fd_sc_hd__inv_2 _08162_ (.A(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__a211o_1 _08163_ (.A1(_02202_),
    .A2(_02209_),
    .B1(_02224_),
    .C1(_02228_),
    .X(_02231_));
 sky130_fd_sc_hd__nand2_2 _08164_ (.A(_02229_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_1 _08165_ (.A(_02225_),
    .B(_02227_),
    .Y(_02233_));
 sky130_fd_sc_hd__xor2_1 _08166_ (.A(_02221_),
    .B(_02222_),
    .X(_02234_));
 sky130_fd_sc_hd__a22o_1 _08167_ (.A1(net866),
    .A2(net2678),
    .B1(_02212_),
    .B2(_02213_),
    .X(_02235_));
 sky130_fd_sc_hd__and4_1 _08168_ (.A(net884),
    .B(net1603),
    .C(net1164),
    .D(net2678),
    .X(_02236_));
 sky130_fd_sc_hd__nand3_1 _08169_ (.A(_02214_),
    .B(_02235_),
    .C(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__a22oi_1 _08170_ (.A1(net977),
    .A2(net734),
    .B1(net1176),
    .B2(net2247),
    .Y(_02238_));
 sky130_fd_sc_hd__and4_1 _08171_ (.A(net2247),
    .B(net977),
    .C(net734),
    .D(net1176),
    .X(_02239_));
 sky130_fd_sc_hd__nor2_1 _08172_ (.A(_02238_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _08173_ (.A(net1160),
    .B(net2674),
    .Y(_02241_));
 sky130_fd_sc_hd__xnor2_1 _08174_ (.A(_02240_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21o_1 _08175_ (.A1(_02214_),
    .A2(_02235_),
    .B1(_02236_),
    .X(_02243_));
 sky130_fd_sc_hd__and3_1 _08176_ (.A(_02237_),
    .B(_02242_),
    .C(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__a21boi_1 _08177_ (.A1(_02242_),
    .A2(_02243_),
    .B1_N(_02237_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2b_1 _08178_ (.A_N(_02245_),
    .B(_02234_),
    .Y(_02246_));
 sky130_fd_sc_hd__o21ba_1 _08179_ (.A1(_02238_),
    .A2(_02241_),
    .B1_N(_02239_),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _08180_ (.A(net1385),
    .B(net2682),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _08181_ (.A(_02247_),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__xnor2_1 _08182_ (.A(_02247_),
    .B(_02248_),
    .Y(_02250_));
 sky130_fd_sc_hd__xor2_1 _08183_ (.A(_02234_),
    .B(_02245_),
    .X(_02251_));
 sky130_fd_sc_hd__o21ai_1 _08184_ (.A1(_02250_),
    .A2(_02251_),
    .B1(_02246_),
    .Y(_02252_));
 sky130_fd_sc_hd__and2_1 _08185_ (.A(_02233_),
    .B(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__xor2_1 _08186_ (.A(_02233_),
    .B(_02252_),
    .X(_02254_));
 sky130_fd_sc_hd__and2_1 _08187_ (.A(_02249_),
    .B(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__or2_2 _08188_ (.A(_02253_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__o21ba_1 _08189_ (.A1(_02253_),
    .A2(_02255_),
    .B1_N(_02232_),
    .X(_02257_));
 sky130_fd_sc_hd__o21ba_1 _08190_ (.A1(_02230_),
    .A2(_02257_),
    .B1_N(_02208_),
    .X(_02258_));
 sky130_fd_sc_hd__xnor2_1 _08191_ (.A(_02249_),
    .B(_02254_),
    .Y(_02259_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(_02250_),
    .B(_02251_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21oi_1 _08193_ (.A1(_02237_),
    .A2(_02243_),
    .B1(_02242_),
    .Y(_02261_));
 sky130_fd_sc_hd__a22o_1 _08194_ (.A1(net866),
    .A2(net734),
    .B1(net1176),
    .B2(net2256),
    .X(_02262_));
 sky130_fd_sc_hd__nand4_2 _08195_ (.A(net977),
    .B(net866),
    .C(net734),
    .D(net1176),
    .Y(_02263_));
 sky130_fd_sc_hd__and2_1 _08196_ (.A(net2247),
    .B(net2674),
    .X(_02264_));
 sky130_fd_sc_hd__a21o_1 _08197_ (.A1(_02262_),
    .A2(_02263_),
    .B1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__nand3_1 _08198_ (.A(_02262_),
    .B(_02263_),
    .C(_02264_),
    .Y(_02266_));
 sky130_fd_sc_hd__a22oi_1 _08199_ (.A1(net1603),
    .A2(net1164),
    .B1(net2678),
    .B2(net1756),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _08200_ (.A(_02236_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand3_1 _08201_ (.A(_02265_),
    .B(_02266_),
    .C(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__or3_1 _08202_ (.A(_02244_),
    .B(_02261_),
    .C(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__a21bo_1 _08203_ (.A1(_02262_),
    .A2(_02264_),
    .B1_N(_02263_),
    .X(_02271_));
 sky130_fd_sc_hd__a21oi_1 _08204_ (.A1(net537),
    .A2(net2682),
    .B1(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__and3_1 _08205_ (.A(net537),
    .B(net2682),
    .C(_02271_),
    .X(_02273_));
 sky130_fd_sc_hd__nor2_1 _08206_ (.A(_02272_),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(net1385),
    .B(net905),
    .Y(_02275_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_02274_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__o21ai_1 _08209_ (.A1(_02244_),
    .A2(_02261_),
    .B1(_02269_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand3_1 _08210_ (.A(_02270_),
    .B(_02276_),
    .C(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _08211_ (.A(_02270_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2b_1 _08212_ (.A_N(_02260_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__a31o_1 _08213_ (.A1(net1385),
    .A2(net905),
    .A3(_02274_),
    .B1(_02273_),
    .X(_02281_));
 sky130_fd_sc_hd__xnor2_1 _08214_ (.A(_02260_),
    .B(_02279_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand2_1 _08215_ (.A(_02281_),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__a21oi_1 _08216_ (.A1(_02280_),
    .A2(_02283_),
    .B1(_02259_),
    .Y(_02284_));
 sky130_fd_sc_hd__nand3_1 _08217_ (.A(_02259_),
    .B(_02280_),
    .C(_02283_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2b_1 _08218_ (.A_N(_02284_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__xnor2_1 _08219_ (.A(_02281_),
    .B(_02282_),
    .Y(_02287_));
 sky130_fd_sc_hd__a21o_1 _08220_ (.A1(_02270_),
    .A2(_02277_),
    .B1(_02276_),
    .X(_02288_));
 sky130_fd_sc_hd__a21o_1 _08221_ (.A1(_02265_),
    .A2(_02266_),
    .B1(_02268_),
    .X(_02289_));
 sky130_fd_sc_hd__nand2_1 _08222_ (.A(net1603),
    .B(net2678),
    .Y(_02290_));
 sky130_fd_sc_hd__a22oi_1 _08223_ (.A1(net1756),
    .A2(net734),
    .B1(net1176),
    .B2(net866),
    .Y(_02291_));
 sky130_fd_sc_hd__a22o_1 _08224_ (.A1(net884),
    .A2(net734),
    .B1(net1176),
    .B2(net866),
    .X(_02292_));
 sky130_fd_sc_hd__and4_1 _08225_ (.A(net866),
    .B(net884),
    .C(net734),
    .D(net1176),
    .X(_02293_));
 sky130_fd_sc_hd__and4b_1 _08226_ (.A_N(_02293_),
    .B(net2674),
    .C(net977),
    .D(_02292_),
    .X(_02294_));
 sky130_fd_sc_hd__o2bb2a_1 _08227_ (.A1_N(net977),
    .A2_N(net2674),
    .B1(_02291_),
    .B2(_02293_),
    .X(_02295_));
 sky130_fd_sc_hd__nor3_1 _08228_ (.A(_02290_),
    .B(_02294_),
    .C(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand3_1 _08229_ (.A(_02269_),
    .B(_02289_),
    .C(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_1 _08230_ (.A(net537),
    .B(net905),
    .Y(_02298_));
 sky130_fd_sc_hd__a31o_1 _08231_ (.A1(net977),
    .A2(net2674),
    .A3(_02292_),
    .B1(_02293_),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_1 _08232_ (.A(net1160),
    .B(net2682),
    .Y(_02300_));
 sky130_fd_sc_hd__and3_1 _08233_ (.A(net1160),
    .B(net2682),
    .C(_02299_),
    .X(_02301_));
 sky130_fd_sc_hd__xnor2_1 _08234_ (.A(_02299_),
    .B(_02300_),
    .Y(_02302_));
 sky130_fd_sc_hd__and3_1 _08235_ (.A(net537),
    .B(net905),
    .C(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__xnor2_1 _08236_ (.A(_02298_),
    .B(_02302_),
    .Y(_02304_));
 sky130_fd_sc_hd__a21o_1 _08237_ (.A1(_02269_),
    .A2(_02289_),
    .B1(_02296_),
    .X(_02305_));
 sky130_fd_sc_hd__nand3_1 _08238_ (.A(_02297_),
    .B(_02304_),
    .C(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand2_1 _08239_ (.A(_02297_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand3_1 _08240_ (.A(_02278_),
    .B(_02288_),
    .C(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a21o_1 _08241_ (.A1(_02278_),
    .A2(_02288_),
    .B1(_02307_),
    .X(_02309_));
 sky130_fd_sc_hd__o211ai_2 _08242_ (.A1(_02301_),
    .A2(_02303_),
    .B1(_02308_),
    .C1(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand2_1 _08243_ (.A(_02308_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__and2b_1 _08244_ (.A_N(_02287_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__xnor2_1 _08245_ (.A(_02287_),
    .B(_02311_),
    .Y(_02313_));
 sky130_fd_sc_hd__a211o_1 _08246_ (.A1(_02308_),
    .A2(_02309_),
    .B1(_02301_),
    .C1(_02303_),
    .X(_02314_));
 sky130_fd_sc_hd__a21o_1 _08247_ (.A1(_02297_),
    .A2(_02305_),
    .B1(_02304_),
    .X(_02315_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(net1160),
    .B(net905),
    .Y(_02316_));
 sky130_fd_sc_hd__and4_1 _08249_ (.A(net884),
    .B(net1603),
    .C(net734),
    .D(net1176),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(net1792),
    .B(net2674),
    .Y(_02318_));
 sky130_fd_sc_hd__a22oi_2 _08251_ (.A1(net1603),
    .A2(net734),
    .B1(net1176),
    .B2(net884),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _08252_ (.A(_02317_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__o21bai_2 _08253_ (.A1(_02318_),
    .A2(_02319_),
    .B1_N(_02317_),
    .Y(_02321_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(net2247),
    .B(net2682),
    .Y(_02322_));
 sky130_fd_sc_hd__and3_1 _08255_ (.A(net2247),
    .B(net2682),
    .C(_02321_),
    .X(_02323_));
 sky130_fd_sc_hd__xnor2_2 _08256_ (.A(_02321_),
    .B(_02322_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _08257_ (.A(_02316_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__o21a_1 _08258_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02290_),
    .X(_02326_));
 sky130_fd_sc_hd__nor2_1 _08259_ (.A(_02296_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__and2_1 _08260_ (.A(_02325_),
    .B(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__and3_1 _08261_ (.A(_02306_),
    .B(_02315_),
    .C(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a31oi_2 _08262_ (.A1(net1160),
    .A2(net3671),
    .A3(_02324_),
    .B1(_02323_),
    .Y(_02330_));
 sky130_fd_sc_hd__a21oi_1 _08263_ (.A1(_02306_),
    .A2(_02315_),
    .B1(_02328_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor3_1 _08264_ (.A(_02329_),
    .B(_02330_),
    .C(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__or3_1 _08265_ (.A(_02329_),
    .B(_02330_),
    .C(_02331_),
    .X(_02333_));
 sky130_fd_sc_hd__o211a_1 _08266_ (.A1(_02329_),
    .A2(_02332_),
    .B1(_02310_),
    .C1(_02314_),
    .X(_02334_));
 sky130_fd_sc_hd__a211o_1 _08267_ (.A1(_02310_),
    .A2(_02314_),
    .B1(_02329_),
    .C1(_02332_),
    .X(_02335_));
 sky130_fd_sc_hd__o21ai_1 _08268_ (.A1(_02329_),
    .A2(_02331_),
    .B1(_02330_),
    .Y(_02336_));
 sky130_fd_sc_hd__xnor2_1 _08269_ (.A(_02325_),
    .B(_02327_),
    .Y(_02337_));
 sky130_fd_sc_hd__xnor2_1 _08270_ (.A(_02318_),
    .B(_02320_),
    .Y(_02338_));
 sky130_fd_sc_hd__and4_1 _08271_ (.A(net884),
    .B(net1603),
    .C(net1176),
    .D(net2674),
    .X(_02339_));
 sky130_fd_sc_hd__inv_2 _08272_ (.A(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__a21oi_1 _08273_ (.A1(net977),
    .A2(net2682),
    .B1(_02339_),
    .Y(_02341_));
 sky130_fd_sc_hd__and3_1 _08274_ (.A(net977),
    .B(net2682),
    .C(_02339_),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _08275_ (.A(_02341_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _08276_ (.A(net2247),
    .B(net905),
    .Y(_02344_));
 sky130_fd_sc_hd__xnor2_1 _08277_ (.A(_02343_),
    .B(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_1 _08278_ (.A(_02338_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _08279_ (.A(_02337_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__a31o_1 _08280_ (.A1(net2247),
    .A2(net905),
    .A3(_02343_),
    .B1(_02342_),
    .X(_02348_));
 sky130_fd_sc_hd__xor2_1 _08281_ (.A(_02337_),
    .B(_02346_),
    .X(_02349_));
 sky130_fd_sc_hd__and2_1 _08282_ (.A(_02348_),
    .B(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__o211a_1 _08283_ (.A1(_02347_),
    .A2(_02350_),
    .B1(_02333_),
    .C1(_02336_),
    .X(_02351_));
 sky130_fd_sc_hd__a211o_1 _08284_ (.A1(_02333_),
    .A2(_02336_),
    .B1(_02347_),
    .C1(_02350_),
    .X(_02352_));
 sky130_fd_sc_hd__nand2b_1 _08285_ (.A_N(_02351_),
    .B(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__xnor2_1 _08286_ (.A(_02348_),
    .B(_02349_),
    .Y(_02354_));
 sky130_fd_sc_hd__xor2_1 _08287_ (.A(_02338_),
    .B(_02345_),
    .X(_02355_));
 sky130_fd_sc_hd__and4_1 _08288_ (.A(net977),
    .B(net866),
    .C(net2682),
    .D(net905),
    .X(_02356_));
 sky130_fd_sc_hd__inv_2 _08289_ (.A(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__a22o_1 _08290_ (.A1(net1603),
    .A2(net1176),
    .B1(net2674),
    .B2(net884),
    .X(_02358_));
 sky130_fd_sc_hd__a22o_1 _08291_ (.A1(net866),
    .A2(net2682),
    .B1(net905),
    .B2(net977),
    .X(_02359_));
 sky130_fd_sc_hd__or4bb_1 _08292_ (.A(_02339_),
    .B(_02356_),
    .C_N(_02358_),
    .D_N(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _08293_ (.A(_02357_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_02355_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _08295_ (.A(_02355_),
    .B(_02361_),
    .Y(_02363_));
 sky130_fd_sc_hd__a22o_1 _08296_ (.A1(_02340_),
    .A2(_02358_),
    .B1(_02359_),
    .B2(_02357_),
    .X(_02364_));
 sky130_fd_sc_hd__and4_1 _08297_ (.A(net866),
    .B(net884),
    .C(net2682),
    .D(net905),
    .X(_02365_));
 sky130_fd_sc_hd__a22o_1 _08298_ (.A1(net884),
    .A2(net2682),
    .B1(net905),
    .B2(net866),
    .X(_02366_));
 sky130_fd_sc_hd__inv_2 _08299_ (.A(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__and4b_1 _08300_ (.A_N(_02365_),
    .B(_02366_),
    .C(net1603),
    .D(net2674),
    .X(_02368_));
 sky130_fd_sc_hd__or2_1 _08301_ (.A(_02365_),
    .B(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__and3_1 _08302_ (.A(_02360_),
    .B(_02364_),
    .C(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__o2bb2a_1 _08303_ (.A1_N(net1603),
    .A2_N(net2674),
    .B1(_02365_),
    .B2(_02367_),
    .X(_02371_));
 sky130_fd_sc_hd__nor2_1 _08304_ (.A(_02368_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__and4_1 _08305_ (.A(net884),
    .B(net1603),
    .C(net2682),
    .D(net905),
    .X(_02373_));
 sky130_fd_sc_hd__and2_1 _08306_ (.A(_02372_),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__a21oi_1 _08307_ (.A1(_02360_),
    .A2(_02364_),
    .B1(_02369_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _08308_ (.A(_02370_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__and2_1 _08309_ (.A(_02374_),
    .B(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__nor2_1 _08310_ (.A(_02370_),
    .B(_02377_),
    .Y(_02378_));
 sky130_fd_sc_hd__o21bai_1 _08311_ (.A1(_02370_),
    .A2(_02377_),
    .B1_N(_02363_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_1 _08312_ (.A1(_02362_),
    .A2(_02379_),
    .B1(_02354_),
    .Y(_02380_));
 sky130_fd_sc_hd__a21o_1 _08313_ (.A1(_02352_),
    .A2(_02380_),
    .B1(_02351_),
    .X(_02381_));
 sky130_fd_sc_hd__a21o_1 _08314_ (.A1(_02335_),
    .A2(_02381_),
    .B1(_02334_),
    .X(_02382_));
 sky130_fd_sc_hd__a21o_1 _08315_ (.A1(_02313_),
    .A2(_02382_),
    .B1(_02312_),
    .X(_02383_));
 sky130_fd_sc_hd__a21o_2 _08316_ (.A1(_02285_),
    .A2(_02383_),
    .B1(_02284_),
    .X(_02384_));
 sky130_fd_sc_hd__xnor2_4 _08317_ (.A(_02232_),
    .B(_02256_),
    .Y(_02385_));
 sky130_fd_sc_hd__xnor2_4 _08318_ (.A(_02208_),
    .B(_02230_),
    .Y(_02386_));
 sky130_fd_sc_hd__a31o_1 _08319_ (.A1(_02384_),
    .A2(_02385_),
    .A3(_02386_),
    .B1(_02258_),
    .X(_02387_));
 sky130_fd_sc_hd__a21oi_2 _08320_ (.A1(_02207_),
    .A2(_02387_),
    .B1(_02205_),
    .Y(_02388_));
 sky130_fd_sc_hd__o21a_1 _08321_ (.A1(_02180_),
    .A2(_02388_),
    .B1(_02178_),
    .X(_02389_));
 sky130_fd_sc_hd__and2b_1 _08322_ (.A_N(_02389_),
    .B(_02153_),
    .X(_02390_));
 sky130_fd_sc_hd__xnor2_2 _08323_ (.A(_02153_),
    .B(_02389_),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(net702),
    .B(net728),
    .Y(_02392_));
 sky130_fd_sc_hd__and4_1 _08325_ (.A(net702),
    .B(net1122),
    .C(net1999),
    .D(net728),
    .X(_02393_));
 sky130_fd_sc_hd__a22o_1 _08326_ (.A1(net1122),
    .A2(net1999),
    .B1(net728),
    .B2(net702),
    .X(_02394_));
 sky130_fd_sc_hd__nand2b_1 _08327_ (.A_N(_02393_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_1 _08328_ (.A(net1452),
    .B(net1942),
    .Y(_02396_));
 sky130_fd_sc_hd__a31o_1 _08329_ (.A1(net1452),
    .A2(net1942),
    .A3(_02394_),
    .B1(_02393_),
    .X(_02397_));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(net702),
    .B(net1999),
    .Y(_02398_));
 sky130_fd_sc_hd__nand2_1 _08331_ (.A(net1452),
    .B(net728),
    .Y(_02399_));
 sky130_fd_sc_hd__xor2_1 _08332_ (.A(_02398_),
    .B(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(_02397_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__or2_1 _08334_ (.A(_02397_),
    .B(_02400_),
    .X(_02402_));
 sky130_fd_sc_hd__nand2_1 _08335_ (.A(_02401_),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__xnor2_1 _08336_ (.A(_02395_),
    .B(_02396_),
    .Y(_02404_));
 sky130_fd_sc_hd__and4_1 _08337_ (.A(net1122),
    .B(net923),
    .C(net1999),
    .D(net728),
    .X(_02405_));
 sky130_fd_sc_hd__inv_2 _08338_ (.A(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__a22o_1 _08339_ (.A1(net923),
    .A2(net1999),
    .B1(net2162),
    .B2(net1122),
    .X(_02407_));
 sky130_fd_sc_hd__and4_1 _08340_ (.A(net702),
    .B(net1942),
    .C(_02406_),
    .D(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__nor2_1 _08341_ (.A(_02405_),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__or2_1 _08342_ (.A(_02404_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_1 _08343_ (.A(_02404_),
    .B(_02409_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _08344_ (.A(_02410_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__a22oi_1 _08345_ (.A1(net702),
    .A2(net1942),
    .B1(_02406_),
    .B2(_02407_),
    .Y(_02413_));
 sky130_fd_sc_hd__or2_1 _08346_ (.A(_02408_),
    .B(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__nand4_2 _08347_ (.A(net923),
    .B(net103),
    .C(net1999),
    .D(net728),
    .Y(_02415_));
 sky130_fd_sc_hd__a22o_1 _08348_ (.A1(net103),
    .A2(net1999),
    .B1(net728),
    .B2(net923),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_1 _08349_ (.A(_02415_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_1 _08350_ (.A(net1122),
    .B(net1942),
    .Y(_02418_));
 sky130_fd_sc_hd__o21ai_2 _08351_ (.A1(_02417_),
    .A2(_02418_),
    .B1(_02415_),
    .Y(_02419_));
 sky130_fd_sc_hd__and2b_1 _08352_ (.A_N(_02414_),
    .B(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__xnor2_1 _08353_ (.A(_02414_),
    .B(_02419_),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(net1452),
    .B(net851),
    .Y(_02422_));
 sky130_fd_sc_hd__a31oi_1 _08355_ (.A1(net1452),
    .A2(net851),
    .A3(_02421_),
    .B1(_02420_),
    .Y(_02423_));
 sky130_fd_sc_hd__or2_1 _08356_ (.A(_02412_),
    .B(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__nor2_1 _08357_ (.A(_02403_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__and2_1 _08358_ (.A(net1452),
    .B(net1999),
    .X(_02426_));
 sky130_fd_sc_hd__nand2_1 _08359_ (.A(_02392_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__o21ai_1 _08360_ (.A1(_02403_),
    .A2(_02410_),
    .B1(_02401_),
    .Y(_02428_));
 sky130_fd_sc_hd__xnor2_1 _08361_ (.A(_02427_),
    .B(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_1 _08362_ (.A(_02425_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _08363_ (.A(_02412_),
    .B(_02423_),
    .Y(_02431_));
 sky130_fd_sc_hd__and2_1 _08364_ (.A(_02424_),
    .B(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__xnor2_1 _08365_ (.A(_02421_),
    .B(_02422_),
    .Y(_02433_));
 sky130_fd_sc_hd__xnor2_1 _08366_ (.A(_02417_),
    .B(_02418_),
    .Y(_02434_));
 sky130_fd_sc_hd__and4_1 _08367_ (.A(net103),
    .B(net104),
    .C(net1999),
    .D(net728),
    .X(_02435_));
 sky130_fd_sc_hd__a22o_1 _08368_ (.A1(net104),
    .A2(net1999),
    .B1(net728),
    .B2(net103),
    .X(_02436_));
 sky130_fd_sc_hd__nand2b_1 _08369_ (.A_N(_02435_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__nand2_1 _08370_ (.A(net923),
    .B(net1942),
    .Y(_02438_));
 sky130_fd_sc_hd__a31o_1 _08371_ (.A1(net923),
    .A2(net1942),
    .A3(_02436_),
    .B1(_02435_),
    .X(_02439_));
 sky130_fd_sc_hd__nand2b_1 _08372_ (.A_N(_02434_),
    .B(_02439_),
    .Y(_02440_));
 sky130_fd_sc_hd__xor2_1 _08373_ (.A(_02434_),
    .B(_02439_),
    .X(_02441_));
 sky130_fd_sc_hd__a22oi_2 _08374_ (.A1(net702),
    .A2(net851),
    .B1(net974),
    .B2(net1452),
    .Y(_02442_));
 sky130_fd_sc_hd__and4_1 _08375_ (.A(net1452),
    .B(net702),
    .C(net851),
    .D(net974),
    .X(_02443_));
 sky130_fd_sc_hd__nor2_1 _08376_ (.A(_02442_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__o31a_1 _08377_ (.A1(_02441_),
    .A2(_02442_),
    .A3(_02443_),
    .B1(_02440_),
    .X(_02445_));
 sky130_fd_sc_hd__and2b_1 _08378_ (.A_N(_02445_),
    .B(_02433_),
    .X(_02446_));
 sky130_fd_sc_hd__xnor2_1 _08379_ (.A(_02433_),
    .B(_02445_),
    .Y(_02447_));
 sky130_fd_sc_hd__a21oi_1 _08380_ (.A1(_02443_),
    .A2(_02447_),
    .B1(_02446_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2b_1 _08381_ (.A_N(_02448_),
    .B(_02432_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _08382_ (.A(_02410_),
    .B(_02424_),
    .Y(_02450_));
 sky130_fd_sc_hd__xor2_1 _08383_ (.A(_02403_),
    .B(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__nor2_1 _08384_ (.A(_02449_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__or2_1 _08385_ (.A(_02449_),
    .B(_02451_),
    .X(_02453_));
 sky130_fd_sc_hd__and2_1 _08386_ (.A(_02449_),
    .B(_02451_),
    .X(_02454_));
 sky130_fd_sc_hd__nor2_1 _08387_ (.A(_02452_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2b_1 _08388_ (.A_N(_02432_),
    .B(_02448_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_02449_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__xnor2_1 _08390_ (.A(_02443_),
    .B(_02447_),
    .Y(_02458_));
 sky130_fd_sc_hd__xnor2_1 _08391_ (.A(_02441_),
    .B(_02444_),
    .Y(_02459_));
 sky130_fd_sc_hd__xnor2_2 _08392_ (.A(_02437_),
    .B(_02438_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand4_2 _08393_ (.A(net104),
    .B(net105),
    .C(net1999),
    .D(net728),
    .Y(_02461_));
 sky130_fd_sc_hd__a22o_1 _08394_ (.A1(net105),
    .A2(net1999),
    .B1(net728),
    .B2(net104),
    .X(_02462_));
 sky130_fd_sc_hd__nand4_2 _08395_ (.A(net103),
    .B(net1942),
    .C(_02461_),
    .D(_02462_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _08396_ (.A(_02461_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__and2b_1 _08397_ (.A_N(_02460_),
    .B(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__a22o_1 _08398_ (.A1(net1122),
    .A2(net851),
    .B1(net974),
    .B2(net702),
    .X(_02466_));
 sky130_fd_sc_hd__and4_1 _08399_ (.A(net702),
    .B(net1122),
    .C(net851),
    .D(net974),
    .X(_02467_));
 sky130_fd_sc_hd__nand4_1 _08400_ (.A(net1531),
    .B(net1122),
    .C(net851),
    .D(net974),
    .Y(_02468_));
 sky130_fd_sc_hd__a22oi_1 _08401_ (.A1(net1452),
    .A2(net947),
    .B1(_02466_),
    .B2(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__and4_1 _08402_ (.A(net1452),
    .B(net947),
    .C(_02466_),
    .D(_02468_),
    .X(_02470_));
 sky130_fd_sc_hd__or2_1 _08403_ (.A(_02469_),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__xor2_2 _08404_ (.A(_02460_),
    .B(_02464_),
    .X(_02472_));
 sky130_fd_sc_hd__nor2_1 _08405_ (.A(_02471_),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__o21a_1 _08406_ (.A1(_02465_),
    .A2(_02473_),
    .B1(_02459_),
    .X(_02474_));
 sky130_fd_sc_hd__o21ai_1 _08407_ (.A1(_02465_),
    .A2(_02473_),
    .B1(_02459_),
    .Y(_02475_));
 sky130_fd_sc_hd__or3_1 _08408_ (.A(_02459_),
    .B(_02465_),
    .C(_02473_),
    .X(_02476_));
 sky130_fd_sc_hd__o211a_1 _08409_ (.A1(_02467_),
    .A2(_02470_),
    .B1(_02475_),
    .C1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__nor2_1 _08410_ (.A(_02474_),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__or2_1 _08411_ (.A(_02458_),
    .B(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__nor2_1 _08412_ (.A(_02457_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__and2_1 _08413_ (.A(_02457_),
    .B(_02479_),
    .X(_02481_));
 sky130_fd_sc_hd__nor2_2 _08414_ (.A(_02480_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _08415_ (.A(_02458_),
    .B(_02478_),
    .Y(_02483_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_02479_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__a211oi_1 _08417_ (.A1(_02475_),
    .A2(_02476_),
    .B1(_02467_),
    .C1(_02470_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_2 _08418_ (.A(_02477_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__xor2_2 _08419_ (.A(_02471_),
    .B(_02472_),
    .X(_02487_));
 sky130_fd_sc_hd__a22o_1 _08420_ (.A1(net103),
    .A2(net1942),
    .B1(_02461_),
    .B2(_02462_),
    .X(_02488_));
 sky130_fd_sc_hd__nand4_1 _08421_ (.A(net105),
    .B(net1648),
    .C(net1999),
    .D(net728),
    .Y(_02489_));
 sky130_fd_sc_hd__and2_1 _08422_ (.A(net104),
    .B(net1942),
    .X(_02490_));
 sky130_fd_sc_hd__a22o_1 _08423_ (.A1(net1648),
    .A2(net1999),
    .B1(net728),
    .B2(net105),
    .X(_02491_));
 sky130_fd_sc_hd__nand3_1 _08424_ (.A(_02489_),
    .B(_02490_),
    .C(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__a21bo_1 _08425_ (.A1(_02490_),
    .A2(_02491_),
    .B1_N(_02489_),
    .X(_02493_));
 sky130_fd_sc_hd__nand3_1 _08426_ (.A(_02463_),
    .B(_02488_),
    .C(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__and4_1 _08427_ (.A(net1122),
    .B(net923),
    .C(net2127),
    .D(net2118),
    .X(_02495_));
 sky130_fd_sc_hd__a22o_1 _08428_ (.A1(net923),
    .A2(net2127),
    .B1(net2118),
    .B2(net2656),
    .X(_02496_));
 sky130_fd_sc_hd__and2b_1 _08429_ (.A_N(_02495_),
    .B(_02496_),
    .X(_02497_));
 sky130_fd_sc_hd__nand2_1 _08430_ (.A(net702),
    .B(net947),
    .Y(_02498_));
 sky130_fd_sc_hd__xnor2_1 _08431_ (.A(_02497_),
    .B(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__a21o_1 _08432_ (.A1(_02463_),
    .A2(_02488_),
    .B1(_02493_),
    .X(_02500_));
 sky130_fd_sc_hd__and3_1 _08433_ (.A(_02494_),
    .B(_02499_),
    .C(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__a31o_1 _08434_ (.A1(_02463_),
    .A2(_02488_),
    .A3(_02493_),
    .B1(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(_02487_),
    .B(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__a31oi_4 _08436_ (.A1(net1531),
    .A2(net947),
    .A3(_02496_),
    .B1(_02495_),
    .Y(_02504_));
 sky130_fd_sc_hd__nor2_1 _08437_ (.A(_02487_),
    .B(_02502_),
    .Y(_02505_));
 sky130_fd_sc_hd__xor2_1 _08438_ (.A(_02487_),
    .B(_02502_),
    .X(_02506_));
 sky130_fd_sc_hd__o21ai_4 _08439_ (.A1(_02504_),
    .A2(_02505_),
    .B1(_02503_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _08440_ (.A(_02486_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__xnor2_4 _08441_ (.A(_02486_),
    .B(_02507_),
    .Y(_02509_));
 sky130_fd_sc_hd__xnor2_1 _08442_ (.A(_02504_),
    .B(_02506_),
    .Y(_02510_));
 sky130_fd_sc_hd__a21oi_1 _08443_ (.A1(_02494_),
    .A2(_02500_),
    .B1(_02499_),
    .Y(_02511_));
 sky130_fd_sc_hd__a21o_1 _08444_ (.A1(_02489_),
    .A2(_02491_),
    .B1(_02490_),
    .X(_02512_));
 sky130_fd_sc_hd__and4_1 _08445_ (.A(net105),
    .B(net1648),
    .C(net728),
    .D(net1942),
    .X(_02513_));
 sky130_fd_sc_hd__inv_2 _08446_ (.A(_02513_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand3_1 _08447_ (.A(_02492_),
    .B(_02512_),
    .C(_02513_),
    .Y(_02515_));
 sky130_fd_sc_hd__and4_1 _08448_ (.A(net2355),
    .B(net103),
    .C(net851),
    .D(net974),
    .X(_02516_));
 sky130_fd_sc_hd__a22o_1 _08449_ (.A1(net103),
    .A2(net2127),
    .B1(net2118),
    .B2(net2355),
    .X(_02517_));
 sky130_fd_sc_hd__and2b_1 _08450_ (.A_N(_02516_),
    .B(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(net1122),
    .B(net947),
    .Y(_02519_));
 sky130_fd_sc_hd__xnor2_1 _08452_ (.A(_02518_),
    .B(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21o_1 _08453_ (.A1(_02492_),
    .A2(_02512_),
    .B1(_02513_),
    .X(_02521_));
 sky130_fd_sc_hd__nand3_1 _08454_ (.A(_02515_),
    .B(_02520_),
    .C(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__a21bo_1 _08455_ (.A1(_02520_),
    .A2(_02521_),
    .B1_N(_02515_),
    .X(_02523_));
 sky130_fd_sc_hd__nor3b_1 _08456_ (.A(_02501_),
    .B(_02511_),
    .C_N(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__a31oi_2 _08457_ (.A1(net1122),
    .A2(net947),
    .A3(_02517_),
    .B1(_02516_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _08458_ (.A(net1452),
    .B(net2045),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _08459_ (.A(_02525_),
    .B(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__xnor2_1 _08460_ (.A(_02525_),
    .B(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21ba_1 _08461_ (.A1(_02501_),
    .A2(_02511_),
    .B1_N(_02523_),
    .X(_02529_));
 sky130_fd_sc_hd__nor3_1 _08462_ (.A(_02524_),
    .B(_02528_),
    .C(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _08463_ (.A(_02524_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__and2b_1 _08464_ (.A_N(_02531_),
    .B(_02510_),
    .X(_02532_));
 sky130_fd_sc_hd__xnor2_1 _08465_ (.A(_02510_),
    .B(_02531_),
    .Y(_02533_));
 sky130_fd_sc_hd__and2_1 _08466_ (.A(_02527_),
    .B(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__or2_2 _08467_ (.A(_02532_),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__o21bai_1 _08468_ (.A1(_02532_),
    .A2(_02534_),
    .B1_N(_02509_),
    .Y(_02536_));
 sky130_fd_sc_hd__a21oi_1 _08469_ (.A1(_02508_),
    .A2(_02536_),
    .B1(_02484_),
    .Y(_02537_));
 sky130_fd_sc_hd__xor2_2 _08470_ (.A(_02484_),
    .B(_02508_),
    .X(_02538_));
 sky130_fd_sc_hd__xnor2_4 _08471_ (.A(_02509_),
    .B(_02535_),
    .Y(_02539_));
 sky130_fd_sc_hd__xnor2_1 _08472_ (.A(_02527_),
    .B(_02533_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21a_1 _08473_ (.A1(_02524_),
    .A2(_02529_),
    .B1(_02528_),
    .X(_02541_));
 sky130_fd_sc_hd__or2_1 _08474_ (.A(_02530_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__a21o_1 _08475_ (.A1(_02515_),
    .A2(_02521_),
    .B1(_02520_),
    .X(_02543_));
 sky130_fd_sc_hd__and4_1 _08476_ (.A(net103),
    .B(net104),
    .C(net851),
    .D(net974),
    .X(_02544_));
 sky130_fd_sc_hd__nand4_2 _08477_ (.A(net103),
    .B(net104),
    .C(net851),
    .D(net974),
    .Y(_02545_));
 sky130_fd_sc_hd__a22o_1 _08478_ (.A1(net104),
    .A2(net851),
    .B1(net974),
    .B2(net103),
    .X(_02546_));
 sky130_fd_sc_hd__and4_1 _08479_ (.A(net923),
    .B(net947),
    .C(_02545_),
    .D(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__nand4_2 _08480_ (.A(net923),
    .B(net947),
    .C(_02545_),
    .D(_02546_),
    .Y(_02548_));
 sky130_fd_sc_hd__a22o_1 _08481_ (.A1(net923),
    .A2(net947),
    .B1(_02545_),
    .B2(_02546_),
    .X(_02549_));
 sky130_fd_sc_hd__a22o_1 _08482_ (.A1(net1648),
    .A2(net728),
    .B1(net1942),
    .B2(net105),
    .X(_02550_));
 sky130_fd_sc_hd__nand4_2 _08483_ (.A(_02514_),
    .B(_02548_),
    .C(_02549_),
    .D(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand3b_1 _08484_ (.A_N(_02551_),
    .B(_02543_),
    .C(_02522_),
    .Y(_02552_));
 sky130_fd_sc_hd__o211a_1 _08485_ (.A1(_02544_),
    .A2(_02547_),
    .B1(net702),
    .C1(net2045),
    .X(_02553_));
 sky130_fd_sc_hd__a211oi_1 _08486_ (.A1(net702),
    .A2(net2045),
    .B1(_02544_),
    .C1(_02547_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _08487_ (.A(_02553_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(net1452),
    .B(net959),
    .Y(_02556_));
 sky130_fd_sc_hd__xnor2_1 _08489_ (.A(_02555_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__a21bo_1 _08490_ (.A1(_02522_),
    .A2(_02543_),
    .B1_N(_02551_),
    .X(_02558_));
 sky130_fd_sc_hd__nand3_1 _08491_ (.A(_02552_),
    .B(_02557_),
    .C(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _08492_ (.A(_02552_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand2b_1 _08493_ (.A_N(_02542_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__a31o_1 _08494_ (.A1(net1452),
    .A2(net959),
    .A3(_02555_),
    .B1(_02553_),
    .X(_02562_));
 sky130_fd_sc_hd__xnor2_1 _08495_ (.A(_02542_),
    .B(_02560_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(_02562_),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__nand3_2 _08497_ (.A(_02540_),
    .B(_02561_),
    .C(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__inv_2 _08498_ (.A(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _08499_ (.A1(_02561_),
    .A2(_02564_),
    .B1(_02540_),
    .Y(_02567_));
 sky130_fd_sc_hd__xnor2_1 _08500_ (.A(_02562_),
    .B(_02563_),
    .Y(_02568_));
 sky130_fd_sc_hd__a21o_1 _08501_ (.A1(_02552_),
    .A2(_02558_),
    .B1(_02557_),
    .X(_02569_));
 sky130_fd_sc_hd__a22o_1 _08502_ (.A1(_02548_),
    .A2(_02549_),
    .B1(_02550_),
    .B2(_02514_),
    .X(_02570_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(net1648),
    .B(net1942),
    .Y(_02571_));
 sky130_fd_sc_hd__and4_1 _08504_ (.A(net104),
    .B(net105),
    .C(net851),
    .D(net974),
    .X(_02572_));
 sky130_fd_sc_hd__a22oi_1 _08505_ (.A1(net105),
    .A2(net851),
    .B1(net974),
    .B2(net104),
    .Y(_02573_));
 sky130_fd_sc_hd__a22o_1 _08506_ (.A1(net105),
    .A2(net851),
    .B1(net974),
    .B2(net104),
    .X(_02574_));
 sky130_fd_sc_hd__and4b_1 _08507_ (.A_N(_02572_),
    .B(_02574_),
    .C(net103),
    .D(net947),
    .X(_02575_));
 sky130_fd_sc_hd__o2bb2a_1 _08508_ (.A1_N(net103),
    .A2_N(net947),
    .B1(_02572_),
    .B2(_02573_),
    .X(_02576_));
 sky130_fd_sc_hd__nor3_2 _08509_ (.A(_02571_),
    .B(_02575_),
    .C(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__and3_1 _08510_ (.A(_02551_),
    .B(_02570_),
    .C(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__nand3_1 _08511_ (.A(_02551_),
    .B(_02570_),
    .C(_02577_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(net702),
    .B(net959),
    .Y(_02580_));
 sky130_fd_sc_hd__a31o_1 _08513_ (.A1(net103),
    .A2(net947),
    .A3(_02574_),
    .B1(_02572_),
    .X(_02581_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(net1122),
    .B(net2045),
    .Y(_02582_));
 sky130_fd_sc_hd__xnor2_1 _08515_ (.A(_02581_),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__and3_1 _08516_ (.A(net702),
    .B(net959),
    .C(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__xnor2_1 _08517_ (.A(_02580_),
    .B(_02583_),
    .Y(_02585_));
 sky130_fd_sc_hd__a21o_1 _08518_ (.A1(_02551_),
    .A2(_02570_),
    .B1(_02577_),
    .X(_02586_));
 sky130_fd_sc_hd__and3_1 _08519_ (.A(_02579_),
    .B(_02585_),
    .C(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__o211ai_2 _08520_ (.A1(_02578_),
    .A2(_02587_),
    .B1(_02559_),
    .C1(_02569_),
    .Y(_02588_));
 sky130_fd_sc_hd__a31o_1 _08521_ (.A1(net1122),
    .A2(net2045),
    .A3(_02581_),
    .B1(_02584_),
    .X(_02589_));
 sky130_fd_sc_hd__a211o_1 _08522_ (.A1(_02559_),
    .A2(_02569_),
    .B1(_02578_),
    .C1(_02587_),
    .X(_02590_));
 sky130_fd_sc_hd__nand3_1 _08523_ (.A(_02588_),
    .B(_02589_),
    .C(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _08524_ (.A(_02588_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__and2b_1 _08525_ (.A_N(_02568_),
    .B(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__a21o_1 _08526_ (.A1(_02588_),
    .A2(_02590_),
    .B1(_02589_),
    .X(_02594_));
 sky130_fd_sc_hd__a21oi_1 _08527_ (.A1(_02579_),
    .A2(_02586_),
    .B1(_02585_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _08528_ (.A(net1122),
    .B(net959),
    .Y(_02596_));
 sky130_fd_sc_hd__and4_1 _08529_ (.A(net105),
    .B(net1648),
    .C(net851),
    .D(net2118),
    .X(_02597_));
 sky130_fd_sc_hd__nand2_1 _08530_ (.A(net104),
    .B(net2193),
    .Y(_02598_));
 sky130_fd_sc_hd__a22oi_1 _08531_ (.A1(net1648),
    .A2(net2127),
    .B1(net974),
    .B2(net1333),
    .Y(_02599_));
 sky130_fd_sc_hd__nor2_1 _08532_ (.A(_02597_),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__o21bai_1 _08533_ (.A1(_02598_),
    .A2(_02599_),
    .B1_N(_02597_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(net923),
    .B(net2045),
    .Y(_02602_));
 sky130_fd_sc_hd__and3_1 _08535_ (.A(net923),
    .B(net2045),
    .C(_02601_),
    .X(_02603_));
 sky130_fd_sc_hd__xnor2_1 _08536_ (.A(_02601_),
    .B(_02602_),
    .Y(_02604_));
 sky130_fd_sc_hd__xnor2_1 _08537_ (.A(_02596_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__o21a_1 _08538_ (.A1(_02575_),
    .A2(_02576_),
    .B1(_02571_),
    .X(_02606_));
 sky130_fd_sc_hd__nor2_1 _08539_ (.A(_02577_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_1 _08540_ (.A(_02605_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__nor3_2 _08541_ (.A(_02587_),
    .B(_02595_),
    .C(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__a31o_1 _08542_ (.A1(net1122),
    .A2(net959),
    .A3(_02604_),
    .B1(_02603_),
    .X(_02610_));
 sky130_fd_sc_hd__inv_2 _08543_ (.A(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__o21a_1 _08544_ (.A1(_02587_),
    .A2(_02595_),
    .B1(_02608_),
    .X(_02612_));
 sky130_fd_sc_hd__nor3_1 _08545_ (.A(_02609_),
    .B(_02611_),
    .C(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__or3_1 _08546_ (.A(_02609_),
    .B(_02611_),
    .C(_02612_),
    .X(_02614_));
 sky130_fd_sc_hd__o211a_1 _08547_ (.A1(_02609_),
    .A2(_02613_),
    .B1(_02591_),
    .C1(_02594_),
    .X(_02615_));
 sky130_fd_sc_hd__a211o_1 _08548_ (.A1(_02591_),
    .A2(_02594_),
    .B1(_02609_),
    .C1(_02613_),
    .X(_02616_));
 sky130_fd_sc_hd__o21ai_1 _08549_ (.A1(_02609_),
    .A2(_02612_),
    .B1(_02611_),
    .Y(_02617_));
 sky130_fd_sc_hd__xnor2_1 _08550_ (.A(_02605_),
    .B(_02607_),
    .Y(_02618_));
 sky130_fd_sc_hd__and4_1 _08551_ (.A(net105),
    .B(net1648),
    .C(net974),
    .D(net2193),
    .X(_02619_));
 sky130_fd_sc_hd__inv_2 _08552_ (.A(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__a21oi_1 _08553_ (.A1(net103),
    .A2(net2045),
    .B1(_02619_),
    .Y(_02621_));
 sky130_fd_sc_hd__and3_1 _08554_ (.A(net1365),
    .B(net2045),
    .C(_02619_),
    .X(_02622_));
 sky130_fd_sc_hd__and4bb_1 _08555_ (.A_N(_02621_),
    .B_N(_02622_),
    .C(net923),
    .D(net959),
    .X(_02623_));
 sky130_fd_sc_hd__o2bb2a_1 _08556_ (.A1_N(net923),
    .A2_N(net959),
    .B1(_02621_),
    .B2(_02622_),
    .X(_02624_));
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(_02623_),
    .B(_02624_),
    .Y(_02625_));
 sky130_fd_sc_hd__xnor2_1 _08558_ (.A(_02598_),
    .B(_02600_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _08559_ (.A(_02625_),
    .B(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__nor2_1 _08560_ (.A(_02618_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__or2_1 _08561_ (.A(_02622_),
    .B(_02623_),
    .X(_02629_));
 sky130_fd_sc_hd__xor2_1 _08562_ (.A(_02618_),
    .B(_02627_),
    .X(_02630_));
 sky130_fd_sc_hd__and2_1 _08563_ (.A(_02629_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__o211a_1 _08564_ (.A1(_02628_),
    .A2(_02631_),
    .B1(_02614_),
    .C1(_02617_),
    .X(_02632_));
 sky130_fd_sc_hd__a211o_1 _08565_ (.A1(_02614_),
    .A2(_02617_),
    .B1(_02628_),
    .C1(_02631_),
    .X(_02633_));
 sky130_fd_sc_hd__nand2b_1 _08566_ (.A_N(_02632_),
    .B(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__xnor2_1 _08567_ (.A(_02629_),
    .B(_02630_),
    .Y(_02635_));
 sky130_fd_sc_hd__xor2_1 _08568_ (.A(_02625_),
    .B(_02626_),
    .X(_02636_));
 sky130_fd_sc_hd__and4_1 _08569_ (.A(net103),
    .B(net104),
    .C(net2045),
    .D(net959),
    .X(_02637_));
 sky130_fd_sc_hd__inv_2 _08570_ (.A(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__a22o_1 _08571_ (.A1(net1648),
    .A2(net974),
    .B1(net947),
    .B2(net105),
    .X(_02639_));
 sky130_fd_sc_hd__a22o_1 _08572_ (.A1(net104),
    .A2(net2045),
    .B1(net959),
    .B2(net1365),
    .X(_02640_));
 sky130_fd_sc_hd__and4_1 _08573_ (.A(_02620_),
    .B(_02638_),
    .C(_02639_),
    .D(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__or4bb_1 _08574_ (.A(_02619_),
    .B(_02637_),
    .C_N(_02639_),
    .D_N(_02640_),
    .X(_02642_));
 sky130_fd_sc_hd__o21ai_2 _08575_ (.A1(_02637_),
    .A2(_02641_),
    .B1(_02636_),
    .Y(_02643_));
 sky130_fd_sc_hd__or3_1 _08576_ (.A(_02636_),
    .B(_02637_),
    .C(_02641_),
    .X(_02644_));
 sky130_fd_sc_hd__a22o_1 _08577_ (.A1(_02620_),
    .A2(_02639_),
    .B1(_02640_),
    .B2(_02638_),
    .X(_02645_));
 sky130_fd_sc_hd__and4_1 _08578_ (.A(net104),
    .B(net105),
    .C(net2045),
    .D(net959),
    .X(_02646_));
 sky130_fd_sc_hd__a22o_1 _08579_ (.A1(net105),
    .A2(net2045),
    .B1(net959),
    .B2(net104),
    .X(_02647_));
 sky130_fd_sc_hd__inv_2 _08580_ (.A(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__and4b_1 _08581_ (.A_N(_02646_),
    .B(_02647_),
    .C(net1648),
    .D(net947),
    .X(_02649_));
 sky130_fd_sc_hd__or2_1 _08582_ (.A(_02646_),
    .B(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__and3_1 _08583_ (.A(_02642_),
    .B(_02645_),
    .C(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__o2bb2a_1 _08584_ (.A1_N(net1648),
    .A2_N(net947),
    .B1(_02646_),
    .B2(_02648_),
    .X(_02652_));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(_02649_),
    .B(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__and4_1 _08586_ (.A(net105),
    .B(net1648),
    .C(net2045),
    .D(net959),
    .X(_02654_));
 sky130_fd_sc_hd__and2_1 _08587_ (.A(_02653_),
    .B(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__a21oi_1 _08588_ (.A1(_02642_),
    .A2(_02645_),
    .B1(_02650_),
    .Y(_02656_));
 sky130_fd_sc_hd__nor2_1 _08589_ (.A(_02651_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__and2_1 _08590_ (.A(_02655_),
    .B(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__o211ai_2 _08591_ (.A1(_02651_),
    .A2(_02658_),
    .B1(_02643_),
    .C1(_02644_),
    .Y(_02659_));
 sky130_fd_sc_hd__a21oi_2 _08592_ (.A1(_02643_),
    .A2(_02659_),
    .B1(_02635_),
    .Y(_02660_));
 sky130_fd_sc_hd__a21o_1 _08593_ (.A1(_02633_),
    .A2(_02660_),
    .B1(_02632_),
    .X(_02661_));
 sky130_fd_sc_hd__a21o_1 _08594_ (.A1(_02616_),
    .A2(_02661_),
    .B1(_02615_),
    .X(_02662_));
 sky130_fd_sc_hd__xnor2_1 _08595_ (.A(_02568_),
    .B(_02592_),
    .Y(_02663_));
 sky130_fd_sc_hd__and2_1 _08596_ (.A(_02662_),
    .B(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__nor2_1 _08597_ (.A(_02593_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__a211o_1 _08598_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_02567_),
    .C1(_02593_),
    .X(_02666_));
 sky130_fd_sc_hd__and2_2 _08599_ (.A(_02565_),
    .B(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__a41o_2 _08600_ (.A1(_02538_),
    .A2(_02539_),
    .A3(_02565_),
    .A4(_02666_),
    .B1(_02537_),
    .X(_02668_));
 sky130_fd_sc_hd__a21oi_1 _08601_ (.A1(_02482_),
    .A2(_02668_),
    .B1(_02480_),
    .Y(_02669_));
 sky130_fd_sc_hd__o21a_1 _08602_ (.A1(_02454_),
    .A2(_02669_),
    .B1(_02453_),
    .X(_02670_));
 sky130_fd_sc_hd__nor2_1 _08603_ (.A(_02430_),
    .B(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__xor2_1 _08604_ (.A(_02430_),
    .B(_02670_),
    .X(_02672_));
 sky130_fd_sc_hd__and2_1 _08605_ (.A(net1514),
    .B(net1917),
    .X(_02673_));
 sky130_fd_sc_hd__a21o_1 _08606_ (.A1(net2209),
    .A2(net163),
    .B1(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__and3_1 _08607_ (.A(net2209),
    .B(net163),
    .C(_02673_),
    .X(_02675_));
 sky130_fd_sc_hd__inv_2 _08608_ (.A(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(_02674_),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(net1500),
    .B(net2123),
    .Y(_02678_));
 sky130_fd_sc_hd__xnor2_1 _08611_ (.A(_02677_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__and4_1 _08612_ (.A(net2209),
    .B(net2179),
    .C(net163),
    .D(net1917),
    .X(_02680_));
 sky130_fd_sc_hd__inv_2 _08613_ (.A(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__a22o_1 _08614_ (.A1(net2179),
    .A2(net163),
    .B1(net1917),
    .B2(net2209),
    .X(_02682_));
 sky130_fd_sc_hd__and4_1 _08615_ (.A(net1514),
    .B(net2123),
    .C(_02681_),
    .D(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__nor2_1 _08616_ (.A(_02680_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__nor2_1 _08617_ (.A(_02679_),
    .B(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__xnor2_1 _08618_ (.A(_02679_),
    .B(_02684_),
    .Y(_02686_));
 sky130_fd_sc_hd__and4_1 _08619_ (.A(net2179),
    .B(net941),
    .C(net163),
    .D(net1917),
    .X(_02687_));
 sky130_fd_sc_hd__inv_2 _08620_ (.A(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__a22o_1 _08621_ (.A1(net941),
    .A2(net163),
    .B1(net1917),
    .B2(net2179),
    .X(_02689_));
 sky130_fd_sc_hd__and4_1 _08622_ (.A(net2209),
    .B(net2123),
    .C(_02688_),
    .D(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__nor2_1 _08623_ (.A(_02687_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__nand2_1 _08624_ (.A(net1500),
    .B(net2091),
    .Y(_02692_));
 sky130_fd_sc_hd__a22oi_1 _08625_ (.A1(net1514),
    .A2(net2123),
    .B1(_02681_),
    .B2(_02682_),
    .Y(_02693_));
 sky130_fd_sc_hd__or2_1 _08626_ (.A(_02683_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__xnor2_1 _08627_ (.A(_02691_),
    .B(_02692_),
    .Y(_02695_));
 sky130_fd_sc_hd__o32a_1 _08628_ (.A1(_02683_),
    .A2(_02693_),
    .A3(_02695_),
    .B1(_02691_),
    .B2(_02692_),
    .X(_02696_));
 sky130_fd_sc_hd__nor2_1 _08629_ (.A(_02686_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__a31o_1 _08630_ (.A1(net1500),
    .A2(net2123),
    .A3(_02674_),
    .B1(_02675_),
    .X(_02698_));
 sky130_fd_sc_hd__a22oi_1 _08631_ (.A1(net1514),
    .A2(net163),
    .B1(net1917),
    .B2(net1500),
    .Y(_02699_));
 sky130_fd_sc_hd__and4_1 _08632_ (.A(net1500),
    .B(net1514),
    .C(net163),
    .D(net1917),
    .X(_02700_));
 sky130_fd_sc_hd__nor2_1 _08633_ (.A(_02699_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__and2_1 _08634_ (.A(_02698_),
    .B(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__nor2_1 _08635_ (.A(_02698_),
    .B(_02701_),
    .Y(_02703_));
 sky130_fd_sc_hd__nor2_1 _08636_ (.A(_02702_),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_1 _08637_ (.A(_02697_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xnor2_1 _08638_ (.A(_02694_),
    .B(_02695_),
    .Y(_02706_));
 sky130_fd_sc_hd__a22oi_1 _08639_ (.A1(net2209),
    .A2(net2123),
    .B1(_02688_),
    .B2(_02689_),
    .Y(_02707_));
 sky130_fd_sc_hd__nor2_1 _08640_ (.A(_02690_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__a22oi_1 _08641_ (.A1(net956),
    .A2(net163),
    .B1(net1917),
    .B2(net941),
    .Y(_02709_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(net956),
    .A2(net163),
    .B1(net1917),
    .B2(net941),
    .X(_02710_));
 sky130_fd_sc_hd__and4_1 _08643_ (.A(net2399),
    .B(net956),
    .C(net163),
    .D(net1917),
    .X(_02711_));
 sky130_fd_sc_hd__o2bb2a_1 _08644_ (.A1_N(net2179),
    .A2_N(net2123),
    .B1(_02709_),
    .B2(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__and4b_1 _08645_ (.A_N(_02711_),
    .B(net2123),
    .C(net2179),
    .D(_02710_),
    .X(_02713_));
 sky130_fd_sc_hd__nor2_2 _08646_ (.A(_02712_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__and2_1 _08647_ (.A(net1514),
    .B(net785),
    .X(_02715_));
 sky130_fd_sc_hd__nand3b_2 _08648_ (.A_N(_02715_),
    .B(net893),
    .C(net1500),
    .Y(_02716_));
 sky130_fd_sc_hd__nand4_2 _08649_ (.A(net1500),
    .B(net1514),
    .C(net893),
    .D(net785),
    .Y(_02717_));
 sky130_fd_sc_hd__o211a_1 _08650_ (.A1(_02714_),
    .A2(_02715_),
    .B1(net1500),
    .C1(net893),
    .X(_02718_));
 sky130_fd_sc_hd__nand2_1 _08651_ (.A(_02708_),
    .B(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__xnor2_1 _08652_ (.A(_02708_),
    .B(_02718_),
    .Y(_02720_));
 sky130_fd_sc_hd__a31o_1 _08653_ (.A1(net2179),
    .A2(net2123),
    .A3(_02710_),
    .B1(_02711_),
    .X(_02721_));
 sky130_fd_sc_hd__a21oi_1 _08654_ (.A1(net1514),
    .A2(net2091),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__and3_1 _08655_ (.A(net1514),
    .B(net2091),
    .C(_02721_),
    .X(_02723_));
 sky130_fd_sc_hd__nor2_1 _08656_ (.A(_02722_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _08657_ (.A(net1500),
    .B(net1833),
    .Y(_02725_));
 sky130_fd_sc_hd__xor2_1 _08658_ (.A(_02724_),
    .B(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__or2_1 _08659_ (.A(_02720_),
    .B(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__a21o_1 _08660_ (.A1(_02719_),
    .A2(_02727_),
    .B1(_02706_),
    .X(_02728_));
 sky130_fd_sc_hd__nand3_1 _08661_ (.A(_02706_),
    .B(_02719_),
    .C(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__and2_1 _08662_ (.A(_02728_),
    .B(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__a31o_1 _08663_ (.A1(net1500),
    .A2(net1833),
    .A3(_02724_),
    .B1(_02723_),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__and2_1 _08665_ (.A(_02686_),
    .B(_02696_),
    .X(_02733_));
 sky130_fd_sc_hd__or2_1 _08666_ (.A(_02697_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__a21o_1 _08667_ (.A1(_02728_),
    .A2(_02732_),
    .B1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__xnor2_2 _08668_ (.A(_02730_),
    .B(_02731_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_1 _08669_ (.A(_02720_),
    .B(_02726_),
    .Y(_02737_));
 sky130_fd_sc_hd__and2_2 _08670_ (.A(_02727_),
    .B(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__xnor2_4 _08671_ (.A(_02714_),
    .B(_02716_),
    .Y(_02739_));
 sky130_fd_sc_hd__a22o_1 _08672_ (.A1(net1514),
    .A2(net893),
    .B1(net785),
    .B2(net1500),
    .X(_02740_));
 sky130_fd_sc_hd__nand2_2 _08673_ (.A(_02717_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand4_2 _08674_ (.A(net1514),
    .B(net2209),
    .C(net893),
    .D(net785),
    .Y(_02742_));
 sky130_fd_sc_hd__and2_1 _08675_ (.A(net1500),
    .B(net1725),
    .X(_02743_));
 sky130_fd_sc_hd__a22o_1 _08676_ (.A1(net2209),
    .A2(net893),
    .B1(net785),
    .B2(net1514),
    .X(_02744_));
 sky130_fd_sc_hd__nand3_1 _08677_ (.A(_02742_),
    .B(_02743_),
    .C(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__a21bo_2 _08678_ (.A1(_02743_),
    .A2(_02744_),
    .B1_N(_02742_),
    .X(_02746_));
 sky130_fd_sc_hd__a22oi_2 _08679_ (.A1(net1829),
    .A2(net1353),
    .B1(net1917),
    .B2(net956),
    .Y(_02747_));
 sky130_fd_sc_hd__and4_1 _08680_ (.A(net956),
    .B(net1829),
    .C(net1353),
    .D(net1917),
    .X(_02748_));
 sky130_fd_sc_hd__nor2_2 _08681_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_2 _08682_ (.A(net2399),
    .B(net2123),
    .Y(_02750_));
 sky130_fd_sc_hd__xnor2_4 _08683_ (.A(_02749_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__xnor2_4 _08684_ (.A(_02741_),
    .B(_02746_),
    .Y(_02752_));
 sky130_fd_sc_hd__a32oi_4 _08685_ (.A1(_02717_),
    .A2(_02740_),
    .A3(_02746_),
    .B1(_02751_),
    .B2(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__and2b_1 _08686_ (.A_N(_02753_),
    .B(_02739_),
    .X(_02754_));
 sky130_fd_sc_hd__o21bai_1 _08687_ (.A1(_02747_),
    .A2(_02750_),
    .B1_N(_02748_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(net2209),
    .B(net2091),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_1 _08689_ (.A(_02755_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__and2_1 _08690_ (.A(net1514),
    .B(net1833),
    .X(_02758_));
 sky130_fd_sc_hd__nor2_1 _08691_ (.A(_02757_),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__and2_1 _08692_ (.A(_02757_),
    .B(_02758_),
    .X(_02760_));
 sky130_fd_sc_hd__nor2_2 _08693_ (.A(_02759_),
    .B(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__xnor2_4 _08694_ (.A(_02739_),
    .B(_02753_),
    .Y(_02762_));
 sky130_fd_sc_hd__a21oi_4 _08695_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_02754_),
    .Y(_02763_));
 sky130_fd_sc_hd__and2b_1 _08696_ (.A_N(_02763_),
    .B(_02738_),
    .X(_02764_));
 sky130_fd_sc_hd__a31o_2 _08697_ (.A1(net2209),
    .A2(net2091),
    .A3(_02755_),
    .B1(_02760_),
    .X(_02765_));
 sky130_fd_sc_hd__xnor2_4 _08698_ (.A(_02738_),
    .B(_02763_),
    .Y(_02766_));
 sky130_fd_sc_hd__a21o_1 _08699_ (.A1(_02765_),
    .A2(_02766_),
    .B1(_02764_),
    .X(_02767_));
 sky130_fd_sc_hd__and2b_1 _08700_ (.A_N(_02736_),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__nand2b_1 _08701_ (.A_N(_02767_),
    .B(_02736_),
    .Y(_02769_));
 sky130_fd_sc_hd__xnor2_2 _08702_ (.A(_02736_),
    .B(_02767_),
    .Y(_02770_));
 sky130_fd_sc_hd__xnor2_4 _08703_ (.A(_02765_),
    .B(_02766_),
    .Y(_02771_));
 sky130_fd_sc_hd__xnor2_2 _08704_ (.A(_02761_),
    .B(_02762_),
    .Y(_02772_));
 sky130_fd_sc_hd__xor2_2 _08705_ (.A(_02751_),
    .B(_02752_),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_1 _08706_ (.A1(net1500),
    .A2(net1725),
    .B1(_02742_),
    .B2(_02744_),
    .X(_02774_));
 sky130_fd_sc_hd__nand4_1 _08707_ (.A(net2209),
    .B(net2179),
    .C(net2852),
    .D(net785),
    .Y(_02775_));
 sky130_fd_sc_hd__and2_1 _08708_ (.A(net1514),
    .B(net1725),
    .X(_02776_));
 sky130_fd_sc_hd__a22o_1 _08709_ (.A1(net2179),
    .A2(net2852),
    .B1(net785),
    .B2(net2209),
    .X(_02777_));
 sky130_fd_sc_hd__nand3_1 _08710_ (.A(_02775_),
    .B(_02776_),
    .C(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__a21bo_1 _08711_ (.A1(_02776_),
    .A2(_02777_),
    .B1_N(_02775_),
    .X(_02779_));
 sky130_fd_sc_hd__nand3_1 _08712_ (.A(_02745_),
    .B(_02774_),
    .C(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(net956),
    .B(net2123),
    .Y(_02781_));
 sky130_fd_sc_hd__a22o_1 _08714_ (.A1(net1640),
    .A2(net163),
    .B1(net1917),
    .B2(net1829),
    .X(_02782_));
 sky130_fd_sc_hd__and3_1 _08715_ (.A(net1829),
    .B(net1640),
    .C(net1917),
    .X(_02783_));
 sky130_fd_sc_hd__a21bo_1 _08716_ (.A1(net163),
    .A2(_02783_),
    .B1_N(_02782_),
    .X(_02784_));
 sky130_fd_sc_hd__xor2_1 _08717_ (.A(_02781_),
    .B(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a21o_1 _08718_ (.A1(_02745_),
    .A2(_02774_),
    .B1(_02779_),
    .X(_02786_));
 sky130_fd_sc_hd__nand3_1 _08719_ (.A(_02780_),
    .B(_02785_),
    .C(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__a21bo_1 _08720_ (.A1(_02785_),
    .A2(_02786_),
    .B1_N(_02780_),
    .X(_02788_));
 sky130_fd_sc_hd__and2_1 _08721_ (.A(_02773_),
    .B(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__a32o_1 _08722_ (.A1(net2183),
    .A2(net2123),
    .A3(_02782_),
    .B1(_02783_),
    .B2(net163),
    .X(_02790_));
 sky130_fd_sc_hd__nand2_1 _08723_ (.A(net2179),
    .B(net2091),
    .Y(_02791_));
 sky130_fd_sc_hd__xnor2_1 _08724_ (.A(_02790_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__and3_1 _08725_ (.A(net2209),
    .B(net1833),
    .C(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__a21oi_1 _08726_ (.A1(net2209),
    .A2(net1833),
    .B1(_02792_),
    .Y(_02794_));
 sky130_fd_sc_hd__nor2_1 _08727_ (.A(_02793_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__xor2_2 _08728_ (.A(_02773_),
    .B(_02788_),
    .X(_02796_));
 sky130_fd_sc_hd__a21o_1 _08729_ (.A1(_02795_),
    .A2(_02796_),
    .B1(_02789_),
    .X(_02797_));
 sky130_fd_sc_hd__and2b_1 _08730_ (.A_N(_02772_),
    .B(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__a31o_1 _08731_ (.A1(net2179),
    .A2(net2091),
    .A3(_02790_),
    .B1(_02793_),
    .X(_02799_));
 sky130_fd_sc_hd__xnor2_2 _08732_ (.A(_02772_),
    .B(_02797_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21oi_2 _08733_ (.A1(_02799_),
    .A2(_02800_),
    .B1(_02798_),
    .Y(_02801_));
 sky130_fd_sc_hd__nor2_1 _08734_ (.A(_02771_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__xor2_4 _08735_ (.A(_02771_),
    .B(_02801_),
    .X(_02803_));
 sky130_fd_sc_hd__xnor2_1 _08736_ (.A(_02799_),
    .B(_02800_),
    .Y(_02804_));
 sky130_fd_sc_hd__xor2_2 _08737_ (.A(_02795_),
    .B(_02796_),
    .X(_02805_));
 sky130_fd_sc_hd__a21o_1 _08738_ (.A1(_02780_),
    .A2(_02786_),
    .B1(_02785_),
    .X(_02806_));
 sky130_fd_sc_hd__a21o_1 _08739_ (.A1(_02775_),
    .A2(_02777_),
    .B1(_02776_),
    .X(_02807_));
 sky130_fd_sc_hd__nand4_1 _08740_ (.A(net2179),
    .B(net941),
    .C(net893),
    .D(net785),
    .Y(_02808_));
 sky130_fd_sc_hd__and2_1 _08741_ (.A(net2209),
    .B(net1725),
    .X(_02809_));
 sky130_fd_sc_hd__a22o_1 _08742_ (.A1(net941),
    .A2(net893),
    .B1(net2105),
    .B2(net2179),
    .X(_02810_));
 sky130_fd_sc_hd__nand3_1 _08743_ (.A(_02808_),
    .B(_02809_),
    .C(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__a21bo_1 _08744_ (.A1(_02809_),
    .A2(_02810_),
    .B1_N(_02808_),
    .X(_02812_));
 sky130_fd_sc_hd__nand3_1 _08745_ (.A(_02778_),
    .B(_02807_),
    .C(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__and2_1 _08746_ (.A(net2123),
    .B(_02783_),
    .X(_02814_));
 sky130_fd_sc_hd__a22oi_1 _08747_ (.A1(net1640),
    .A2(net1917),
    .B1(net2123),
    .B2(net1829),
    .Y(_02815_));
 sky130_fd_sc_hd__nor2_1 _08748_ (.A(_02814_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__a21o_1 _08749_ (.A1(_02778_),
    .A2(_02807_),
    .B1(_02812_),
    .X(_02817_));
 sky130_fd_sc_hd__nand3_1 _08750_ (.A(_02813_),
    .B(_02816_),
    .C(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__a21bo_1 _08751_ (.A1(_02816_),
    .A2(_02817_),
    .B1_N(_02813_),
    .X(_02819_));
 sky130_fd_sc_hd__and3_1 _08752_ (.A(_02787_),
    .B(_02806_),
    .C(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__a21oi_1 _08753_ (.A1(net2401),
    .A2(net2091),
    .B1(_02814_),
    .Y(_02821_));
 sky130_fd_sc_hd__and3_1 _08754_ (.A(net2401),
    .B(net2091),
    .C(_02814_),
    .X(_02822_));
 sky130_fd_sc_hd__or2_1 _08755_ (.A(_02821_),
    .B(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(net2179),
    .B(net1833),
    .Y(_02824_));
 sky130_fd_sc_hd__xor2_1 _08757_ (.A(_02823_),
    .B(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__a21o_1 _08758_ (.A1(_02787_),
    .A2(_02806_),
    .B1(_02819_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2b_1 _08759_ (.A_N(_02820_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__a21o_1 _08760_ (.A1(_02825_),
    .A2(_02826_),
    .B1(_02820_),
    .X(_02828_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_02805_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__o21ba_1 _08762_ (.A1(_02821_),
    .A2(_02824_),
    .B1_N(_02822_),
    .X(_02830_));
 sky130_fd_sc_hd__xor2_2 _08763_ (.A(_02805_),
    .B(_02828_),
    .X(_02831_));
 sky130_fd_sc_hd__nand2b_1 _08764_ (.A_N(_02830_),
    .B(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21oi_1 _08765_ (.A1(_02829_),
    .A2(_02832_),
    .B1(_02804_),
    .Y(_02833_));
 sky130_fd_sc_hd__and3_1 _08766_ (.A(_02804_),
    .B(_02829_),
    .C(_02832_),
    .X(_02834_));
 sky130_fd_sc_hd__xnor2_2 _08767_ (.A(_02830_),
    .B(_02831_),
    .Y(_02835_));
 sky130_fd_sc_hd__xnor2_1 _08768_ (.A(_02825_),
    .B(_02827_),
    .Y(_02836_));
 sky130_fd_sc_hd__a21o_1 _08769_ (.A1(_02813_),
    .A2(_02817_),
    .B1(_02816_),
    .X(_02837_));
 sky130_fd_sc_hd__a21o_1 _08770_ (.A1(_02808_),
    .A2(_02810_),
    .B1(_02809_),
    .X(_02838_));
 sky130_fd_sc_hd__nand4_2 _08771_ (.A(net941),
    .B(net956),
    .C(net893),
    .D(net785),
    .Y(_02839_));
 sky130_fd_sc_hd__and2_1 _08772_ (.A(net2179),
    .B(net1725),
    .X(_02840_));
 sky130_fd_sc_hd__a22o_1 _08773_ (.A1(net956),
    .A2(net893),
    .B1(net785),
    .B2(net941),
    .X(_02841_));
 sky130_fd_sc_hd__nand3_1 _08774_ (.A(_02839_),
    .B(_02840_),
    .C(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__a21bo_1 _08775_ (.A1(_02840_),
    .A2(_02841_),
    .B1_N(_02839_),
    .X(_02843_));
 sky130_fd_sc_hd__and3_1 _08776_ (.A(_02811_),
    .B(_02838_),
    .C(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_1 _08777_ (.A(net1640),
    .B(net2123),
    .Y(_02845_));
 sky130_fd_sc_hd__a21oi_1 _08778_ (.A1(_02811_),
    .A2(_02838_),
    .B1(_02843_),
    .Y(_02846_));
 sky130_fd_sc_hd__or3_1 _08779_ (.A(_02844_),
    .B(_02845_),
    .C(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__o21bai_1 _08780_ (.A1(_02845_),
    .A2(_02846_),
    .B1_N(_02844_),
    .Y(_02848_));
 sky130_fd_sc_hd__and3_1 _08781_ (.A(_02818_),
    .B(_02837_),
    .C(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__and4_2 _08782_ (.A(net2401),
    .B(net2185),
    .C(net2091),
    .D(net1833),
    .X(_02850_));
 sky130_fd_sc_hd__a22oi_2 _08783_ (.A1(net2185),
    .A2(net2091),
    .B1(net1833),
    .B2(net2401),
    .Y(_02851_));
 sky130_fd_sc_hd__a21oi_1 _08784_ (.A1(_02818_),
    .A2(_02837_),
    .B1(_02848_),
    .Y(_02852_));
 sky130_fd_sc_hd__or4_1 _08785_ (.A(_02849_),
    .B(_02850_),
    .C(_02851_),
    .D(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__and2b_1 _08786_ (.A_N(_02849_),
    .B(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__and2b_1 _08787_ (.A_N(_02854_),
    .B(_02836_),
    .X(_02855_));
 sky130_fd_sc_hd__xnor2_1 _08788_ (.A(_02836_),
    .B(_02854_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21oi_2 _08789_ (.A1(_02850_),
    .A2(_02856_),
    .B1(_02855_),
    .Y(_02857_));
 sky130_fd_sc_hd__and2b_1 _08790_ (.A_N(_02857_),
    .B(_02835_),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _08791_ (.A(_02850_),
    .B(_02856_),
    .Y(_02859_));
 sky130_fd_sc_hd__o22ai_2 _08792_ (.A1(_02850_),
    .A2(_02851_),
    .B1(_02852_),
    .B2(_02849_),
    .Y(_02860_));
 sky130_fd_sc_hd__o21ai_1 _08793_ (.A1(_02844_),
    .A2(_02846_),
    .B1(_02845_),
    .Y(_02861_));
 sky130_fd_sc_hd__and4_1 _08794_ (.A(net956),
    .B(net1829),
    .C(net893),
    .D(net785),
    .X(_02862_));
 sky130_fd_sc_hd__inv_2 _08795_ (.A(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__a22o_1 _08796_ (.A1(net1829),
    .A2(net893),
    .B1(net785),
    .B2(net956),
    .X(_02864_));
 sky130_fd_sc_hd__and4_1 _08797_ (.A(net941),
    .B(net1725),
    .C(_02863_),
    .D(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__a31o_1 _08798_ (.A1(net941),
    .A2(net1725),
    .A3(_02864_),
    .B1(_02862_),
    .X(_02866_));
 sky130_fd_sc_hd__a21o_1 _08799_ (.A1(_02839_),
    .A2(_02841_),
    .B1(_02840_),
    .X(_02867_));
 sky130_fd_sc_hd__and3_1 _08800_ (.A(_02842_),
    .B(_02866_),
    .C(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__nand3_1 _08801_ (.A(_02847_),
    .B(_02861_),
    .C(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__a22oi_1 _08802_ (.A1(net1829),
    .A2(net2091),
    .B1(net1833),
    .B2(net956),
    .Y(_02870_));
 sky130_fd_sc_hd__and4_1 _08803_ (.A(net2185),
    .B(net1829),
    .C(net2091),
    .D(net1833),
    .X(_02871_));
 sky130_fd_sc_hd__nor2_1 _08804_ (.A(_02870_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__a21o_1 _08805_ (.A1(_02847_),
    .A2(_02861_),
    .B1(_02868_),
    .X(_02873_));
 sky130_fd_sc_hd__nand3_1 _08806_ (.A(_02869_),
    .B(_02872_),
    .C(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__a21bo_1 _08807_ (.A1(_02872_),
    .A2(_02873_),
    .B1_N(_02869_),
    .X(_02875_));
 sky130_fd_sc_hd__nand3_2 _08808_ (.A(_02853_),
    .B(_02860_),
    .C(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__a21o_1 _08809_ (.A1(_02853_),
    .A2(_02860_),
    .B1(_02875_),
    .X(_02877_));
 sky130_fd_sc_hd__nand3_2 _08810_ (.A(_02871_),
    .B(_02876_),
    .C(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(_02876_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__and2b_1 _08812_ (.A_N(_02859_),
    .B(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__nand2b_1 _08813_ (.A_N(_02859_),
    .B(_02879_),
    .Y(_02881_));
 sky130_fd_sc_hd__and3_1 _08814_ (.A(_02859_),
    .B(_02876_),
    .C(_02878_),
    .X(_02882_));
 sky130_fd_sc_hd__nor2_1 _08815_ (.A(_02880_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__a21o_1 _08816_ (.A1(_02876_),
    .A2(_02877_),
    .B1(_02871_),
    .X(_02884_));
 sky130_fd_sc_hd__a21o_1 _08817_ (.A1(_02869_),
    .A2(_02873_),
    .B1(_02872_),
    .X(_02885_));
 sky130_fd_sc_hd__a21oi_1 _08818_ (.A1(_02842_),
    .A2(_02867_),
    .B1(_02866_),
    .Y(_02886_));
 sky130_fd_sc_hd__or2_1 _08819_ (.A(_02868_),
    .B(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__a22oi_1 _08820_ (.A1(net941),
    .A2(net1725),
    .B1(_02863_),
    .B2(_02864_),
    .Y(_02888_));
 sky130_fd_sc_hd__and3_1 _08821_ (.A(net1829),
    .B(net1640),
    .C(net785),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(net956),
    .B(net1725),
    .Y(_02890_));
 sky130_fd_sc_hd__a22o_1 _08823_ (.A1(net1640),
    .A2(net893),
    .B1(net785),
    .B2(net1829),
    .X(_02891_));
 sky130_fd_sc_hd__a21bo_1 _08824_ (.A1(net893),
    .A2(_02889_),
    .B1_N(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__o2bb2a_1 _08825_ (.A1_N(net893),
    .A2_N(_02889_),
    .B1(_02890_),
    .B2(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__nor3_1 _08826_ (.A(_02865_),
    .B(_02888_),
    .C(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__and2b_1 _08827_ (.A_N(_02887_),
    .B(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__a22oi_1 _08828_ (.A1(net1640),
    .A2(net2091),
    .B1(net1833),
    .B2(net1829),
    .Y(_02896_));
 sky130_fd_sc_hd__and4_1 _08829_ (.A(net1829),
    .B(net1640),
    .C(net2091),
    .D(net1833),
    .X(_02897_));
 sky130_fd_sc_hd__nor2_1 _08830_ (.A(_02896_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__xnor2_1 _08831_ (.A(_02887_),
    .B(_02894_),
    .Y(_02899_));
 sky130_fd_sc_hd__a21o_1 _08832_ (.A1(_02898_),
    .A2(_02899_),
    .B1(_02895_),
    .X(_02900_));
 sky130_fd_sc_hd__nand3_1 _08833_ (.A(_02874_),
    .B(_02885_),
    .C(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21o_1 _08834_ (.A1(_02874_),
    .A2(_02885_),
    .B1(_02900_),
    .X(_02902_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_02901_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__a21bo_1 _08836_ (.A1(_02897_),
    .A2(_02902_),
    .B1_N(_02901_),
    .X(_02904_));
 sky130_fd_sc_hd__and3_1 _08837_ (.A(_02878_),
    .B(_02884_),
    .C(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__nand3_1 _08838_ (.A(_02878_),
    .B(_02884_),
    .C(_02904_),
    .Y(_02906_));
 sky130_fd_sc_hd__xnor2_1 _08839_ (.A(_02898_),
    .B(_02899_),
    .Y(_02907_));
 sky130_fd_sc_hd__xor2_1 _08840_ (.A(_02890_),
    .B(_02892_),
    .X(_02908_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(net1725),
    .B(_02889_),
    .Y(_02909_));
 sky130_fd_sc_hd__inv_2 _08842_ (.A(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__and2_1 _08843_ (.A(_02908_),
    .B(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__o21a_1 _08844_ (.A1(_02865_),
    .A2(_02888_),
    .B1(_02893_),
    .X(_02912_));
 sky130_fd_sc_hd__nor2_1 _08845_ (.A(_02894_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_02911_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _08847_ (.A(net1640),
    .B(net1833),
    .Y(_02915_));
 sky130_fd_sc_hd__xor2_1 _08848_ (.A(_02911_),
    .B(_02913_),
    .X(_02916_));
 sky130_fd_sc_hd__nand2b_1 _08849_ (.A_N(_02915_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21oi_2 _08850_ (.A1(_02914_),
    .A2(_02917_),
    .B1(_02907_),
    .Y(_02918_));
 sky130_fd_sc_hd__inv_2 _08851_ (.A(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__xor2_1 _08852_ (.A(_02897_),
    .B(_02903_),
    .X(_02920_));
 sky130_fd_sc_hd__or2_1 _08853_ (.A(_02919_),
    .B(_02920_),
    .X(_02921_));
 sky130_fd_sc_hd__a21oi_2 _08854_ (.A1(_02878_),
    .A2(_02884_),
    .B1(_02904_),
    .Y(_02922_));
 sky130_fd_sc_hd__or3_1 _08855_ (.A(_02905_),
    .B(_02921_),
    .C(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__o31a_2 _08856_ (.A1(_02919_),
    .A2(_02920_),
    .A3(_02922_),
    .B1(_02906_),
    .X(_02924_));
 sky130_fd_sc_hd__o21ai_4 _08857_ (.A1(_02882_),
    .A2(_02924_),
    .B1(_02881_),
    .Y(_02925_));
 sky130_fd_sc_hd__xnor2_2 _08858_ (.A(_02835_),
    .B(_02857_),
    .Y(_02926_));
 sky130_fd_sc_hd__a21o_1 _08859_ (.A1(_02925_),
    .A2(_02926_),
    .B1(_02858_),
    .X(_02927_));
 sky130_fd_sc_hd__nor2_1 _08860_ (.A(_02833_),
    .B(_02834_),
    .Y(_02928_));
 sky130_fd_sc_hd__and2_1 _08861_ (.A(_02926_),
    .B(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__o21ba_1 _08862_ (.A1(_02833_),
    .A2(_02858_),
    .B1_N(_02834_),
    .X(_02930_));
 sky130_fd_sc_hd__a21o_1 _08863_ (.A1(_02925_),
    .A2(_02929_),
    .B1(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__and2_1 _08864_ (.A(_02770_),
    .B(_02803_),
    .X(_02932_));
 sky130_fd_sc_hd__nand3_1 _08865_ (.A(_02925_),
    .B(_02929_),
    .C(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_02930_),
    .B(_02932_),
    .Y(_02934_));
 sky130_fd_sc_hd__a21oi_1 _08867_ (.A1(_02769_),
    .A2(_02802_),
    .B1(_02768_),
    .Y(_02935_));
 sky130_fd_sc_hd__nand3_2 _08868_ (.A(_02933_),
    .B(_02934_),
    .C(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand3_1 _08869_ (.A(_02728_),
    .B(_02732_),
    .C(_02734_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand2_2 _08870_ (.A(_02735_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a31o_1 _08871_ (.A1(_02933_),
    .A2(_02934_),
    .A3(_02935_),
    .B1(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__nor3_1 _08872_ (.A(_02685_),
    .B(_02697_),
    .C(_02704_),
    .Y(_02940_));
 sky130_fd_sc_hd__and2_1 _08873_ (.A(_02685_),
    .B(_02704_),
    .X(_02941_));
 sky130_fd_sc_hd__a211o_1 _08874_ (.A1(_02697_),
    .A2(_02704_),
    .B1(_02940_),
    .C1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__a21o_1 _08875_ (.A1(_02735_),
    .A2(_02939_),
    .B1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__or2_1 _08876_ (.A(_02702_),
    .B(_02941_),
    .X(_02944_));
 sky130_fd_sc_hd__and3b_1 _08877_ (.A_N(_02673_),
    .B(net163),
    .C(net1500),
    .X(_02945_));
 sky130_fd_sc_hd__xnor2_1 _08878_ (.A(_02944_),
    .B(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__a21o_1 _08879_ (.A1(_02705_),
    .A2(_02943_),
    .B1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__nand3_1 _08880_ (.A(_02705_),
    .B(_02943_),
    .C(_02946_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand3_1 _08881_ (.A(_02672_),
    .B(_02947_),
    .C(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__a21o_1 _08882_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02672_),
    .X(_02950_));
 sky130_fd_sc_hd__and3_1 _08883_ (.A(_02391_),
    .B(_02949_),
    .C(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__a21oi_1 _08884_ (.A1(_02949_),
    .A2(_02950_),
    .B1(_02391_),
    .Y(_02952_));
 sky130_fd_sc_hd__xnor2_1 _08885_ (.A(_02455_),
    .B(_02669_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand3_1 _08886_ (.A(_02735_),
    .B(_02939_),
    .C(_02942_),
    .Y(_02954_));
 sky130_fd_sc_hd__and3_1 _08887_ (.A(_02943_),
    .B(_02953_),
    .C(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__xnor2_2 _08888_ (.A(_02180_),
    .B(_02388_),
    .Y(_02956_));
 sky130_fd_sc_hd__a21oi_1 _08889_ (.A1(_02943_),
    .A2(_02954_),
    .B1(_02953_),
    .Y(_02957_));
 sky130_fd_sc_hd__nor3_2 _08890_ (.A(_02955_),
    .B(_02956_),
    .C(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nor2_1 _08891_ (.A(_02955_),
    .B(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__nor3_2 _08892_ (.A(_02951_),
    .B(_02952_),
    .C(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__o21a_1 _08893_ (.A1(_02951_),
    .A2(_02952_),
    .B1(_02959_),
    .X(_02961_));
 sky130_fd_sc_hd__or3_1 _08894_ (.A(_02115_),
    .B(_02960_),
    .C(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o21ai_1 _08895_ (.A1(_02960_),
    .A2(_02961_),
    .B1(_02115_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21a_1 _08896_ (.A1(_02955_),
    .A2(_02957_),
    .B1(_02956_),
    .X(_02964_));
 sky130_fd_sc_hd__xnor2_4 _08897_ (.A(_02482_),
    .B(_02668_),
    .Y(_02965_));
 sky130_fd_sc_hd__xor2_4 _08898_ (.A(_02936_),
    .B(_02938_),
    .X(_02966_));
 sky130_fd_sc_hd__or2_1 _08899_ (.A(_02965_),
    .B(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__xor2_2 _08900_ (.A(_02207_),
    .B(_02387_),
    .X(_02968_));
 sky130_fd_sc_hd__inv_2 _08901_ (.A(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__xnor2_4 _08902_ (.A(_02965_),
    .B(_02966_),
    .Y(_02970_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(_02969_),
    .B(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__a211oi_4 _08904_ (.A1(_02967_),
    .A2(_02971_),
    .B1(_02958_),
    .C1(_02964_),
    .Y(_02972_));
 sky130_fd_sc_hd__xor2_2 _08905_ (.A(_02073_),
    .B(_02074_),
    .X(_02973_));
 sky130_fd_sc_hd__o211a_1 _08906_ (.A1(_02958_),
    .A2(_02964_),
    .B1(_02967_),
    .C1(_02971_),
    .X(_02974_));
 sky130_fd_sc_hd__nor3_2 _08907_ (.A(_02972_),
    .B(_02973_),
    .C(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__or2_1 _08908_ (.A(_02972_),
    .B(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__and3_1 _08909_ (.A(_02962_),
    .B(_02963_),
    .C(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__a21oi_1 _08910_ (.A1(_02962_),
    .A2(_02963_),
    .B1(_02976_),
    .Y(_02978_));
 sky130_fd_sc_hd__nor2_1 _08911_ (.A(_02977_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__xnor2_1 _08912_ (.A(_02087_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__o21a_1 _08913_ (.A1(_02972_),
    .A2(_02974_),
    .B1(_02973_),
    .X(_02981_));
 sky130_fd_sc_hd__xnor2_4 _08914_ (.A(_02969_),
    .B(_02970_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21bo_1 _08915_ (.A1(_02539_),
    .A2(_02667_),
    .B1_N(_02536_),
    .X(_02983_));
 sky130_fd_sc_hd__xor2_2 _08916_ (.A(_02538_),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__a21oi_1 _08917_ (.A1(_02803_),
    .A2(_02931_),
    .B1(_02802_),
    .Y(_02985_));
 sky130_fd_sc_hd__xnor2_2 _08918_ (.A(_02770_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__and2_1 _08919_ (.A(_02984_),
    .B(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__or2_1 _08920_ (.A(_02984_),
    .B(_02986_),
    .X(_02988_));
 sky130_fd_sc_hd__xnor2_2 _08921_ (.A(_02984_),
    .B(_02986_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_2 _08922_ (.A1(_02384_),
    .A2(_02385_),
    .B1(_02257_),
    .Y(_02990_));
 sky130_fd_sc_hd__xnor2_4 _08923_ (.A(_02386_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21oi_2 _08924_ (.A1(_02988_),
    .A2(_02991_),
    .B1(_02987_),
    .Y(_02992_));
 sky130_fd_sc_hd__or2_2 _08925_ (.A(_02982_),
    .B(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__nand2_1 _08926_ (.A(_01461_),
    .B(_01462_),
    .Y(_02994_));
 sky130_fd_sc_hd__and2_1 _08927_ (.A(_01463_),
    .B(_02994_),
    .X(_02995_));
 sky130_fd_sc_hd__xor2_4 _08928_ (.A(_02982_),
    .B(_02992_),
    .X(_02996_));
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(_02995_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__a211o_1 _08930_ (.A1(_02993_),
    .A2(_02997_),
    .B1(_02975_),
    .C1(_02981_),
    .X(_02998_));
 sky130_fd_sc_hd__xor2_2 _08931_ (.A(_02020_),
    .B(_02021_),
    .X(_02999_));
 sky130_fd_sc_hd__o211ai_2 _08932_ (.A1(_02975_),
    .A2(_02981_),
    .B1(_02993_),
    .C1(_02997_),
    .Y(_03000_));
 sky130_fd_sc_hd__and3_1 _08933_ (.A(_02998_),
    .B(_02999_),
    .C(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__a21bo_1 _08934_ (.A1(_02999_),
    .A2(_03000_),
    .B1_N(_02998_),
    .X(_03002_));
 sky130_fd_sc_hd__nand2_1 _08935_ (.A(_02980_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__xor2_1 _08936_ (.A(_02980_),
    .B(_03002_),
    .X(_03004_));
 sky130_fd_sc_hd__xnor2_1 _08937_ (.A(_02022_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__a21oi_1 _08938_ (.A1(_02998_),
    .A2(_03000_),
    .B1(_02999_),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_1 _08939_ (.A(_02995_),
    .B(_02996_),
    .Y(_03007_));
 sky130_fd_sc_hd__xnor2_4 _08940_ (.A(_02989_),
    .B(_02991_),
    .Y(_03008_));
 sky130_fd_sc_hd__xor2_4 _08941_ (.A(_02539_),
    .B(_02667_),
    .X(_03009_));
 sky130_fd_sc_hd__xor2_4 _08942_ (.A(_02803_),
    .B(_02931_),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_03009_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__xnor2_4 _08944_ (.A(_02384_),
    .B(_02385_),
    .Y(_03012_));
 sky130_fd_sc_hd__xnor2_4 _08945_ (.A(_03009_),
    .B(_03010_),
    .Y(_03013_));
 sky130_fd_sc_hd__o21a_2 _08946_ (.A1(_03012_),
    .A2(_03013_),
    .B1(_03011_),
    .X(_03014_));
 sky130_fd_sc_hd__and2b_1 _08947_ (.A_N(_03014_),
    .B(_03008_),
    .X(_03015_));
 sky130_fd_sc_hd__a31o_1 _08948_ (.A1(_00824_),
    .A2(_00855_),
    .A3(_00949_),
    .B1(_00820_),
    .X(_03016_));
 sky130_fd_sc_hd__xor2_2 _08949_ (.A(_00823_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__a21oi_2 _08950_ (.A1(_01081_),
    .A2(_01208_),
    .B1(_01078_),
    .Y(_03018_));
 sky130_fd_sc_hd__xnor2_4 _08951_ (.A(_01080_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_03017_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__xnor2_2 _08953_ (.A(_03017_),
    .B(_03019_),
    .Y(_03021_));
 sky130_fd_sc_hd__xnor2_2 _08954_ (.A(_01304_),
    .B(_01458_),
    .Y(_03022_));
 sky130_fd_sc_hd__xnor2_4 _08955_ (.A(_01303_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__or2_1 _08956_ (.A(_03021_),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__xnor2_2 _08957_ (.A(_03021_),
    .B(_03023_),
    .Y(_03025_));
 sky130_fd_sc_hd__inv_2 _08958_ (.A(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__xnor2_4 _08959_ (.A(_03008_),
    .B(_03014_),
    .Y(_03027_));
 sky130_fd_sc_hd__a21oi_1 _08960_ (.A1(_03026_),
    .A2(_03027_),
    .B1(_03015_),
    .Y(_03028_));
 sky130_fd_sc_hd__or2_1 _08961_ (.A(_03007_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__or3_1 _08962_ (.A(_01802_),
    .B(_01840_),
    .C(_02007_),
    .X(_03030_));
 sky130_fd_sc_hd__and2_1 _08963_ (.A(_02008_),
    .B(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__nor3_1 _08964_ (.A(_01548_),
    .B(_01575_),
    .C(_01734_),
    .Y(_03032_));
 sky130_fd_sc_hd__or2_2 _08965_ (.A(_01735_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__a21o_1 _08966_ (.A1(_03020_),
    .A2(_03024_),
    .B1(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__nand3_1 _08967_ (.A(_03020_),
    .B(_03024_),
    .C(_03033_),
    .Y(_03035_));
 sky130_fd_sc_hd__and2_1 _08968_ (.A(_03034_),
    .B(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_03031_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__xnor2_1 _08970_ (.A(_03031_),
    .B(_03036_),
    .Y(_03038_));
 sky130_fd_sc_hd__xnor2_1 _08971_ (.A(_03007_),
    .B(_03028_),
    .Y(_03039_));
 sky130_fd_sc_hd__or2_1 _08972_ (.A(_03038_),
    .B(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a211oi_2 _08973_ (.A1(_03029_),
    .A2(_03040_),
    .B1(_03001_),
    .C1(_03006_),
    .Y(_03041_));
 sky130_fd_sc_hd__o211a_1 _08974_ (.A1(_03001_),
    .A2(_03006_),
    .B1(_03029_),
    .C1(_03040_),
    .X(_03042_));
 sky130_fd_sc_hd__a211oi_2 _08975_ (.A1(_03034_),
    .A2(_03037_),
    .B1(_03041_),
    .C1(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__nor2_1 _08976_ (.A(_03041_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_03005_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__xor2_1 _08978_ (.A(_03005_),
    .B(_03044_),
    .X(_03046_));
 sky130_fd_sc_hd__o211a_1 _08979_ (.A1(_03041_),
    .A2(_03042_),
    .B1(_03034_),
    .C1(_03037_),
    .X(_03047_));
 sky130_fd_sc_hd__xnor2_1 _08980_ (.A(_03038_),
    .B(_03039_),
    .Y(_03048_));
 sky130_fd_sc_hd__xnor2_1 _08981_ (.A(_03025_),
    .B(_03027_),
    .Y(_03049_));
 sky130_fd_sc_hd__xnor2_4 _08982_ (.A(_03012_),
    .B(_03013_),
    .Y(_03050_));
 sky130_fd_sc_hd__or2_1 _08983_ (.A(_02566_),
    .B(_02567_),
    .X(_03051_));
 sky130_fd_sc_hd__xnor2_2 _08984_ (.A(_02665_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__xnor2_2 _08985_ (.A(_02927_),
    .B(_02928_),
    .Y(_03053_));
 sky130_fd_sc_hd__nor2_1 _08986_ (.A(_03052_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__xor2_2 _08987_ (.A(_02286_),
    .B(_02383_),
    .X(_03055_));
 sky130_fd_sc_hd__inv_2 _08988_ (.A(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__xor2_2 _08989_ (.A(_03052_),
    .B(_03053_),
    .X(_03057_));
 sky130_fd_sc_hd__a21oi_2 _08990_ (.A1(_03056_),
    .A2(_03057_),
    .B1(_03054_),
    .Y(_03058_));
 sky130_fd_sc_hd__xnor2_2 _08991_ (.A(_01331_),
    .B(_01457_),
    .Y(_03059_));
 sky130_fd_sc_hd__xnor2_2 _08992_ (.A(_00824_),
    .B(_00950_),
    .Y(_03060_));
 sky130_fd_sc_hd__xnor2_2 _08993_ (.A(_01081_),
    .B(_01208_),
    .Y(_03061_));
 sky130_fd_sc_hd__inv_2 _08994_ (.A(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_1 _08995_ (.A(_03060_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__xnor2_1 _08996_ (.A(_03060_),
    .B(_03062_),
    .Y(_03064_));
 sky130_fd_sc_hd__or2_1 _08997_ (.A(_03059_),
    .B(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__xor2_1 _08998_ (.A(_03059_),
    .B(_03064_),
    .X(_03066_));
 sky130_fd_sc_hd__xor2_1 _08999_ (.A(_03050_),
    .B(_03058_),
    .X(_03067_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(_03066_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__o21a_1 _09001_ (.A1(_03050_),
    .A2(_03058_),
    .B1(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2b_1 _09002_ (.A_N(_03069_),
    .B(_03049_),
    .Y(_03070_));
 sky130_fd_sc_hd__and3_1 _09003_ (.A(_01842_),
    .B(_01872_),
    .C(_02006_),
    .X(_03071_));
 sky130_fd_sc_hd__or2_1 _09004_ (.A(_02007_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__and3_1 _09005_ (.A(_01577_),
    .B(_01609_),
    .C(_01733_),
    .X(_03073_));
 sky130_fd_sc_hd__or2_1 _09006_ (.A(_01734_),
    .B(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__a21oi_1 _09007_ (.A1(_03063_),
    .A2(_03065_),
    .B1(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__a21o_1 _09008_ (.A1(_03063_),
    .A2(_03065_),
    .B1(_03074_),
    .X(_03076_));
 sky130_fd_sc_hd__and3_1 _09009_ (.A(_03063_),
    .B(_03065_),
    .C(_03074_),
    .X(_03077_));
 sky130_fd_sc_hd__nor2_1 _09010_ (.A(_03075_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__xnor2_1 _09011_ (.A(_03072_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__xnor2_1 _09012_ (.A(_03049_),
    .B(_03069_),
    .Y(_03080_));
 sky130_fd_sc_hd__a21boi_1 _09013_ (.A1(_03079_),
    .A2(_03080_),
    .B1_N(_03070_),
    .Y(_03081_));
 sky130_fd_sc_hd__or2_1 _09014_ (.A(_03048_),
    .B(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__o21a_1 _09015_ (.A1(_03072_),
    .A2(_03077_),
    .B1(_03076_),
    .X(_03083_));
 sky130_fd_sc_hd__xor2_1 _09016_ (.A(_03048_),
    .B(_03081_),
    .X(_03084_));
 sky130_fd_sc_hd__nand2b_1 _09017_ (.A_N(_03083_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__o211a_1 _09018_ (.A1(_03043_),
    .A2(_03047_),
    .B1(_03082_),
    .C1(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__a211o_1 _09019_ (.A1(_03082_),
    .A2(_03085_),
    .B1(_03043_),
    .C1(_03047_),
    .X(_03087_));
 sky130_fd_sc_hd__xnor2_1 _09020_ (.A(_03083_),
    .B(_03084_),
    .Y(_03088_));
 sky130_fd_sc_hd__xnor2_1 _09021_ (.A(_03079_),
    .B(_03080_),
    .Y(_03089_));
 sky130_fd_sc_hd__xnor2_1 _09022_ (.A(_03066_),
    .B(_03067_),
    .Y(_03090_));
 sky130_fd_sc_hd__xnor2_2 _09023_ (.A(_03055_),
    .B(_03057_),
    .Y(_03091_));
 sky130_fd_sc_hd__nor2_1 _09024_ (.A(_02662_),
    .B(_02663_),
    .Y(_03092_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(_02664_),
    .B(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__xor2_2 _09026_ (.A(_02925_),
    .B(_02926_),
    .X(_03094_));
 sky130_fd_sc_hd__and2b_1 _09027_ (.A_N(_03093_),
    .B(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__xnor2_1 _09028_ (.A(_02313_),
    .B(_02382_),
    .Y(_03096_));
 sky130_fd_sc_hd__xor2_1 _09029_ (.A(_03093_),
    .B(_03094_),
    .X(_03097_));
 sky130_fd_sc_hd__nor2_1 _09030_ (.A(_03096_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__nor2_1 _09031_ (.A(_03095_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__and2b_1 _09032_ (.A_N(_03099_),
    .B(_03091_),
    .X(_03100_));
 sky130_fd_sc_hd__xnor2_2 _09033_ (.A(_01358_),
    .B(_01456_),
    .Y(_03101_));
 sky130_fd_sc_hd__xnor2_2 _09034_ (.A(_01109_),
    .B(_01207_),
    .Y(_03102_));
 sky130_fd_sc_hd__nor2_1 _09035_ (.A(_00854_),
    .B(_00856_),
    .Y(_03103_));
 sky130_fd_sc_hd__xnor2_2 _09036_ (.A(_00948_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hd__xor2_2 _09037_ (.A(_03102_),
    .B(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__nand2b_1 _09038_ (.A_N(_03101_),
    .B(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__xnor2_2 _09039_ (.A(_03101_),
    .B(_03105_),
    .Y(_03107_));
 sky130_fd_sc_hd__xnor2_2 _09040_ (.A(_03091_),
    .B(_03099_),
    .Y(_03108_));
 sky130_fd_sc_hd__a21oi_1 _09041_ (.A1(_03107_),
    .A2(_03108_),
    .B1(_03100_),
    .Y(_03109_));
 sky130_fd_sc_hd__nor2_1 _09042_ (.A(_03090_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand3_1 _09043_ (.A(net3460),
    .B(_01901_),
    .C(_02005_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_02006_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__o21a_1 _09045_ (.A1(_03102_),
    .A2(_03104_),
    .B1(_03106_),
    .X(_03113_));
 sky130_fd_sc_hd__or3_1 _09046_ (.A(_01610_),
    .B(_01636_),
    .C(_01732_),
    .X(_03114_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(_01733_),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__xnor2_1 _09048_ (.A(_03113_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__nor2_1 _09049_ (.A(_03112_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__xor2_1 _09050_ (.A(_03112_),
    .B(_03116_),
    .X(_03118_));
 sky130_fd_sc_hd__xor2_1 _09051_ (.A(_03090_),
    .B(_03109_),
    .X(_03119_));
 sky130_fd_sc_hd__a21o_1 _09052_ (.A1(_03118_),
    .A2(_03119_),
    .B1(_03110_),
    .X(_03120_));
 sky130_fd_sc_hd__and2b_1 _09053_ (.A_N(_03089_),
    .B(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o21bai_2 _09054_ (.A1(_03113_),
    .A2(_03115_),
    .B1_N(_03117_),
    .Y(_03122_));
 sky130_fd_sc_hd__xor2_1 _09055_ (.A(_03089_),
    .B(_03120_),
    .X(_03123_));
 sky130_fd_sc_hd__and2b_1 _09056_ (.A_N(_03123_),
    .B(_03122_),
    .X(_03124_));
 sky130_fd_sc_hd__o21ai_1 _09057_ (.A1(_03121_),
    .A2(_03124_),
    .B1(_03088_),
    .Y(_03125_));
 sky130_fd_sc_hd__a21oi_1 _09058_ (.A1(_03087_),
    .A2(_03125_),
    .B1(_03086_),
    .Y(_03126_));
 sky130_fd_sc_hd__and2b_1 _09059_ (.A_N(_03086_),
    .B(_03087_),
    .X(_03127_));
 sky130_fd_sc_hd__or3_1 _09060_ (.A(_03088_),
    .B(_03121_),
    .C(_03124_),
    .X(_03128_));
 sky130_fd_sc_hd__and2_1 _09061_ (.A(_03125_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__xnor2_1 _09062_ (.A(_03122_),
    .B(_03123_),
    .Y(_03130_));
 sky130_fd_sc_hd__xnor2_1 _09063_ (.A(_03118_),
    .B(_03119_),
    .Y(_03131_));
 sky130_fd_sc_hd__xnor2_1 _09064_ (.A(_03107_),
    .B(_03108_),
    .Y(_03132_));
 sky130_fd_sc_hd__xnor2_1 _09065_ (.A(_01384_),
    .B(net3701),
    .Y(_03133_));
 sky130_fd_sc_hd__xor2_2 _09066_ (.A(_00946_),
    .B(_00947_),
    .X(_03134_));
 sky130_fd_sc_hd__inv_2 _09067_ (.A(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__a21oi_1 _09068_ (.A1(_01155_),
    .A2(_01205_),
    .B1(_01133_),
    .Y(_03136_));
 sky130_fd_sc_hd__or2_2 _09069_ (.A(_01206_),
    .B(_03136_),
    .X(_03137_));
 sky130_fd_sc_hd__nor2_1 _09070_ (.A(_03135_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xor2_1 _09071_ (.A(_03134_),
    .B(_03137_),
    .X(_03139_));
 sky130_fd_sc_hd__nor2_1 _09072_ (.A(_03133_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(_03133_),
    .B(_03139_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2b_1 _09074_ (.A_N(_03140_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(_03096_),
    .B(_03097_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2b_2 _09076_ (.A_N(_03098_),
    .B(net2853),
    .Y(_03144_));
 sky130_fd_sc_hd__or2_1 _09077_ (.A(_03142_),
    .B(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__nor2_1 _09078_ (.A(_03132_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand3_1 _09079_ (.A(_01902_),
    .B(_01927_),
    .C(_02004_),
    .Y(_03147_));
 sky130_fd_sc_hd__and2_1 _09080_ (.A(_02005_),
    .B(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__o211a_1 _09081_ (.A1(_01636_),
    .A2(_01637_),
    .B1(_01662_),
    .C1(_01731_),
    .X(_03149_));
 sky130_fd_sc_hd__nor2_1 _09082_ (.A(_01732_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__o21a_1 _09083_ (.A1(_03138_),
    .A2(_03140_),
    .B1(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__nor3_1 _09084_ (.A(_03138_),
    .B(_03140_),
    .C(_03150_),
    .Y(_03152_));
 sky130_fd_sc_hd__nor2_1 _09085_ (.A(_03151_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__xnor2_1 _09086_ (.A(_03148_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__inv_2 _09087_ (.A(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__xor2_1 _09088_ (.A(_03132_),
    .B(_03145_),
    .X(_03156_));
 sky130_fd_sc_hd__a21oi_1 _09089_ (.A1(_03155_),
    .A2(_03156_),
    .B1(_03146_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_1 _09090_ (.A1(_03148_),
    .A2(_03153_),
    .B1(_03151_),
    .X(_03158_));
 sky130_fd_sc_hd__xnor2_1 _09091_ (.A(_03131_),
    .B(_03157_),
    .Y(_03159_));
 sky130_fd_sc_hd__and2b_1 _09092_ (.A_N(_03159_),
    .B(_03158_),
    .X(_03160_));
 sky130_fd_sc_hd__o21ba_1 _09093_ (.A1(_03131_),
    .A2(_03157_),
    .B1_N(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__and2b_1 _09094_ (.A_N(_03161_),
    .B(_03130_),
    .X(_03162_));
 sky130_fd_sc_hd__xor2_1 _09095_ (.A(_03158_),
    .B(_03159_),
    .X(_03163_));
 sky130_fd_sc_hd__xnor2_1 _09096_ (.A(_03154_),
    .B(_03156_),
    .Y(_03164_));
 sky130_fd_sc_hd__a211o_1 _09097_ (.A1(_01662_),
    .A2(_01663_),
    .B1(_01684_),
    .C1(_01730_),
    .X(_03165_));
 sky130_fd_sc_hd__nand2_1 _09098_ (.A(_01731_),
    .B(net2779),
    .Y(_03166_));
 sky130_fd_sc_hd__or3_1 _09099_ (.A(_01928_),
    .B(_01950_),
    .C(_02003_),
    .X(_03167_));
 sky130_fd_sc_hd__and2_1 _09100_ (.A(_02004_),
    .B(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nand2b_1 _09101_ (.A_N(net2780),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__inv_2 _09102_ (.A(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(net3702),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _09104_ (.A(_03142_),
    .B(_03144_),
    .Y(_03172_));
 sky130_fd_sc_hd__and2_1 _09105_ (.A(_03145_),
    .B(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__xnor2_1 _09106_ (.A(net2780),
    .B(_03168_),
    .Y(_03174_));
 sky130_fd_sc_hd__and3_1 _09107_ (.A(_03145_),
    .B(net2855),
    .C(net2781),
    .X(_03175_));
 sky130_fd_sc_hd__nand2_1 _09108_ (.A(_03164_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__a21o_1 _09109_ (.A1(_03171_),
    .A2(_03176_),
    .B1(_03163_),
    .X(_03177_));
 sky130_fd_sc_hd__inv_2 _09110_ (.A(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__xnor2_1 _09111_ (.A(_03130_),
    .B(_03161_),
    .Y(_03179_));
 sky130_fd_sc_hd__a21o_1 _09112_ (.A1(_03178_),
    .A2(_03179_),
    .B1(_03162_),
    .X(_03180_));
 sky130_fd_sc_hd__nand2_1 _09113_ (.A(_03129_),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__a31o_1 _09114_ (.A1(_03127_),
    .A2(_03129_),
    .A3(_03180_),
    .B1(_03126_),
    .X(_03182_));
 sky130_fd_sc_hd__a21oi_1 _09115_ (.A1(_03046_),
    .A2(_03182_),
    .B1(_03045_),
    .Y(_03183_));
 sky130_fd_sc_hd__o2bb2a_1 _09116_ (.A1_N(_02107_),
    .A2_N(_02110_),
    .B1(_02111_),
    .B2(_02106_),
    .X(_03184_));
 sky130_fd_sc_hd__a21o_1 _09117_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02102_),
    .X(_03185_));
 sky130_fd_sc_hd__or3b_1 _09118_ (.A(_03185_),
    .B(_02100_),
    .C_N(_02034_),
    .X(_03186_));
 sky130_fd_sc_hd__xnor2_1 _09119_ (.A(_03184_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__a21oi_1 _09120_ (.A1(_02088_),
    .A2(_02089_),
    .B1(_02061_),
    .Y(_03188_));
 sky130_fd_sc_hd__and3_1 _09121_ (.A(_02092_),
    .B(_02094_),
    .C(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__a21oi_1 _09122_ (.A1(_02052_),
    .A2(_02109_),
    .B1(_02049_),
    .Y(_03190_));
 sky130_fd_sc_hd__xnor2_1 _09123_ (.A(_03189_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_2 _09124_ (.A(_03187_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__a21o_1 _09125_ (.A1(_02135_),
    .A2(_02136_),
    .B1(net3601),
    .X(_03193_));
 sky130_fd_sc_hd__a211oi_4 _09126_ (.A1(_02138_),
    .A2(_02152_),
    .B1(_02390_),
    .C1(net3609),
    .Y(_03194_));
 sky130_fd_sc_hd__o211a_1 _09127_ (.A1(_02673_),
    .A2(_02702_),
    .B1(net1500),
    .C1(net163),
    .X(_03195_));
 sky130_fd_sc_hd__nand2b_1 _09128_ (.A_N(_02428_),
    .B(_02392_),
    .Y(_03196_));
 sky130_fd_sc_hd__a221o_1 _09129_ (.A1(_02425_),
    .A2(_02429_),
    .B1(_03196_),
    .B2(_02426_),
    .C1(_02671_),
    .X(_03197_));
 sky130_fd_sc_hd__xor2_1 _09130_ (.A(_03195_),
    .B(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__xnor2_2 _09131_ (.A(net3610),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__xnor2_1 _09132_ (.A(_03192_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o21ba_1 _09133_ (.A1(_02087_),
    .A2(_02978_),
    .B1_N(_02977_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2b_1 _09134_ (.A_N(_02960_),
    .B(_02962_),
    .Y(_03202_));
 sky130_fd_sc_hd__a31o_1 _09135_ (.A1(_02672_),
    .A2(_02947_),
    .A3(_02948_),
    .B1(_02951_),
    .X(_03203_));
 sky130_fd_sc_hd__a21bo_1 _09136_ (.A1(_02941_),
    .A2(_02945_),
    .B1_N(_02947_),
    .X(_03204_));
 sky130_fd_sc_hd__xor2_2 _09137_ (.A(_03203_),
    .B(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__xnor2_1 _09138_ (.A(_03202_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__xnor2_1 _09139_ (.A(_03201_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__xnor2_1 _09140_ (.A(_03200_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__a21boi_1 _09141_ (.A1(_02022_),
    .A2(_03004_),
    .B1_N(_03003_),
    .Y(_03209_));
 sky130_fd_sc_hd__o21a_2 _09142_ (.A1(_02097_),
    .A2(_02114_),
    .B1(_02113_),
    .X(_03210_));
 sky130_fd_sc_hd__a21o_1 _09143_ (.A1(_02078_),
    .A2(_02079_),
    .B1(_02081_),
    .X(_03211_));
 sky130_fd_sc_hd__xnor2_1 _09144_ (.A(_03210_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__and3_1 _09145_ (.A(_02012_),
    .B(_02027_),
    .C(_02030_),
    .X(_03213_));
 sky130_fd_sc_hd__xnor2_1 _09146_ (.A(_03212_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__a21oi_2 _09147_ (.A1(_02076_),
    .A2(_02077_),
    .B1(_01513_),
    .Y(_03215_));
 sky130_fd_sc_hd__nor2_1 _09148_ (.A(_02084_),
    .B(_02086_),
    .Y(_03216_));
 sky130_fd_sc_hd__xnor2_1 _09149_ (.A(_03215_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__xnor2_2 _09150_ (.A(_03214_),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__xnor2_1 _09151_ (.A(_03209_),
    .B(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__xnor2_1 _09152_ (.A(_03208_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__xnor2_1 _09153_ (.A(_03183_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(net1233),
    .A1(_03221_),
    .S(net37),
    .X(_00544_));
 sky130_fd_sc_hd__or2_1 _09155_ (.A(_03046_),
    .B(_03182_),
    .X(_03222_));
 sky130_fd_sc_hd__a21oi_1 _09156_ (.A1(_03046_),
    .A2(_03182_),
    .B1(net34),
    .Y(_03223_));
 sky130_fd_sc_hd__a22o_1 _09157_ (.A1(net1321),
    .A2(net34),
    .B1(_03222_),
    .B2(_03223_),
    .X(_00543_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(net3461),
    .B(_03181_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _09159_ (.A(net3813),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__o21a_1 _09160_ (.A1(_03127_),
    .A2(_03224_),
    .B1(net37),
    .X(_03226_));
 sky130_fd_sc_hd__a22o_1 _09161_ (.A1(net1325),
    .A2(net34),
    .B1(_03225_),
    .B2(_03226_),
    .X(_00542_));
 sky130_fd_sc_hd__and2_1 _09162_ (.A(net2594),
    .B(net34),
    .X(_03227_));
 sky130_fd_sc_hd__or2_1 _09163_ (.A(_03129_),
    .B(_03180_),
    .X(_03228_));
 sky130_fd_sc_hd__a31o_1 _09164_ (.A1(net37),
    .A2(_03181_),
    .A3(_03228_),
    .B1(net2596),
    .X(_00541_));
 sky130_fd_sc_hd__or2_1 _09165_ (.A(_03178_),
    .B(_03179_),
    .X(_03229_));
 sky130_fd_sc_hd__a21oi_1 _09166_ (.A1(_03178_),
    .A2(_03179_),
    .B1(net34),
    .Y(_03230_));
 sky130_fd_sc_hd__a22o_1 _09167_ (.A1(net1317),
    .A2(net34),
    .B1(_03229_),
    .B2(_03230_),
    .X(_00540_));
 sky130_fd_sc_hd__and3_1 _09168_ (.A(_03163_),
    .B(_03171_),
    .C(_03176_),
    .X(_03231_));
 sky130_fd_sc_hd__nand2_1 _09169_ (.A(net37),
    .B(_03177_),
    .Y(_03232_));
 sky130_fd_sc_hd__a2bb2o_1 _09170_ (.A1_N(_03231_),
    .A2_N(_03232_),
    .B1(net1301),
    .B2(net34),
    .X(_00539_));
 sky130_fd_sc_hd__and2_1 _09171_ (.A(net2570),
    .B(net34),
    .X(_03233_));
 sky130_fd_sc_hd__or2_1 _09172_ (.A(_03164_),
    .B(_03175_),
    .X(_03234_));
 sky130_fd_sc_hd__a21o_1 _09173_ (.A1(_03176_),
    .A2(net2857),
    .B1(_03170_),
    .X(_03235_));
 sky130_fd_sc_hd__a31o_1 _09174_ (.A1(net37),
    .A2(net3703),
    .A3(_03235_),
    .B1(net2572),
    .X(_00538_));
 sky130_fd_sc_hd__or2_1 _09175_ (.A(_03173_),
    .B(net2781),
    .X(_03236_));
 sky130_fd_sc_hd__nor2_1 _09176_ (.A(net34),
    .B(_03175_),
    .Y(_03237_));
 sky130_fd_sc_hd__a22o_1 _09177_ (.A1(net1397),
    .A2(net34),
    .B1(net2782),
    .B2(_03237_),
    .X(_00537_));
 sky130_fd_sc_hd__nand2_4 _09178_ (.A(_00676_),
    .B(net1622),
    .Y(_03238_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(net174),
    .A1(net1452),
    .S(_03238_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(net175),
    .A1(net1533),
    .S(_03238_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(net2286),
    .A1(net2658),
    .S(_03238_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(net1014),
    .A1(net2357),
    .S(_03238_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _09183_ (.A0(net1018),
    .A1(net3075),
    .S(_03238_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(net179),
    .A1(net2977),
    .S(_03238_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(net180),
    .A1(net3031),
    .S(_03238_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(net181),
    .A1(net1648),
    .S(_03238_),
    .X(_00529_));
 sky130_fd_sc_hd__or3b_2 _09187_ (.A(net1341),
    .B(net1545),
    .C_N(net1537),
    .X(_03239_));
 sky130_fd_sc_hd__nor3_1 _09188_ (.A(net2407),
    .B(net1893),
    .C(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__mux2_1 _09189_ (.A0(net1709),
    .A1(net2368),
    .S(net2409),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(net1672),
    .A1(net1875),
    .S(net2409),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _09191_ (.A0(net1887),
    .A1(net2327),
    .S(net2409),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(net2449),
    .A1(net1682),
    .S(net2409),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(net2433),
    .A1(net2033),
    .S(net2409),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(net2189),
    .A1(net2087),
    .S(net2409),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(net2427),
    .A1(net1797),
    .S(net2409),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net896),
    .A1(net1922),
    .S(net2409),
    .X(_00521_));
 sky130_fd_sc_hd__nor3b_1 _09197_ (.A(_03239_),
    .B(net2407),
    .C_N(net1893),
    .Y(_03241_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(net1930),
    .A1(net2368),
    .S(net31),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(net2317),
    .A1(net1875),
    .S(net31),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net1938),
    .A1(net2327),
    .S(net31),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net2477),
    .A1(net1682),
    .S(net31),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(net2483),
    .A1(net2033),
    .S(net31),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(net1717),
    .A1(net2087),
    .S(net31),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(net1713),
    .A1(net1797),
    .S(net31),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(net1926),
    .A1(net1922),
    .S(net31),
    .X(_00513_));
 sky130_fd_sc_hd__nor3b_1 _09206_ (.A(net1865),
    .B(_03239_),
    .C_N(net1599),
    .Y(_03242_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(net1857),
    .A1(net2368),
    .S(net1866),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(net675),
    .A1(net1875),
    .S(net1866),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(net1870),
    .A1(net2327),
    .S(net1866),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(net746),
    .A1(net1682),
    .S(net1866),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(net2074),
    .A1(net2033),
    .S(net1866),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(net1690),
    .A1(net2087),
    .S(net1866),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(net1767),
    .A1(net1797),
    .S(net1866),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(net821),
    .A1(net1922),
    .S(net1866),
    .X(_00505_));
 sky130_fd_sc_hd__and2_2 _09215_ (.A(net2407),
    .B(net1893),
    .X(_03243_));
 sky130_fd_sc_hd__and2b_4 _09216_ (.A_N(_03239_),
    .B(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(net3421),
    .A1(net2368),
    .S(_03244_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(net2277),
    .A1(net1875),
    .S(_03244_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(net3347),
    .A1(net2327),
    .S(_03244_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _09220_ (.A0(net2460),
    .A1(net1682),
    .S(_03244_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(net2465),
    .A1(net2033),
    .S(_03244_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _09222_ (.A0(net3553),
    .A1(net2087),
    .S(_03244_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(net1805),
    .A1(net1797),
    .S(_03244_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _09224_ (.A0(net3640),
    .A1(net1922),
    .S(_03244_),
    .X(_00497_));
 sky130_fd_sc_hd__and2b_4 _09225_ (.A_N(net1341),
    .B(net1545),
    .X(_03245_));
 sky130_fd_sc_hd__and4bb_4 _09226_ (.A_N(net1599),
    .B_N(net1893),
    .C(_03245_),
    .D(net1537),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(net3391),
    .A1(net2368),
    .S(_03246_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _09228_ (.A0(net2028),
    .A1(net1875),
    .S(_03246_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(net3313),
    .A1(net2327),
    .S(_03246_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _09230_ (.A0(net2390),
    .A1(net1682),
    .S(_03246_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(net2395),
    .A1(net2033),
    .S(_03246_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _09232_ (.A0(net3531),
    .A1(net2087),
    .S(_03246_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(net1809),
    .A1(net1797),
    .S(_03246_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _09234_ (.A0(net2379),
    .A1(net1922),
    .S(_03246_),
    .X(_00489_));
 sky130_fd_sc_hd__and3b_4 _09235_ (.A_N(net1599),
    .B(net1893),
    .C(net1537),
    .X(_03247_));
 sky130_fd_sc_hd__nand2_8 _09236_ (.A(_03245_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(net2368),
    .A1(net1837),
    .S(_03248_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _09238_ (.A0(net1875),
    .A1(net1743),
    .S(_03248_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _09239_ (.A0(net2327),
    .A1(net872),
    .S(_03248_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(net1682),
    .A1(net2003),
    .S(_03248_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _09241_ (.A0(net2033),
    .A1(net1668),
    .S(_03248_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _09242_ (.A0(net2087),
    .A1(net2363),
    .S(_03248_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(net1797),
    .A1(net2132),
    .S(_03248_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _09244_ (.A0(net1922),
    .A1(net2239),
    .S(_03248_),
    .X(_00481_));
 sky130_fd_sc_hd__and3b_4 _09245_ (.A_N(net1893),
    .B(net1599),
    .C(net1537),
    .X(_03249_));
 sky130_fd_sc_hd__nand2_4 _09246_ (.A(_03245_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(net2368),
    .A1(net3475),
    .S(_03250_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _09248_ (.A0(net1875),
    .A1(net2282),
    .S(_03250_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(net2327),
    .A1(net3369),
    .S(_03250_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _09250_ (.A0(net1682),
    .A1(net3613),
    .S(_03250_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(net2033),
    .A1(net3619),
    .S(_03250_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _09252_ (.A0(net2087),
    .A1(net2298),
    .S(_03250_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(net1797),
    .A1(net1954),
    .S(_03250_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _09254_ (.A0(net1922),
    .A1(net3150),
    .S(_03250_),
    .X(_00473_));
 sky130_fd_sc_hd__and3_4 _09255_ (.A(net1537),
    .B(net1599),
    .C(net1893),
    .X(_03251_));
 sky130_fd_sc_hd__nand2_8 _09256_ (.A(_03245_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(net2368),
    .A1(net3507),
    .S(_03252_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _09258_ (.A0(net1875),
    .A1(net3050),
    .S(_03252_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(net2327),
    .A1(net3442),
    .S(_03252_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _09260_ (.A0(net1682),
    .A1(net3434),
    .S(_03252_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _09261_ (.A0(net2033),
    .A1(net2876),
    .S(_03252_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _09262_ (.A0(net2087),
    .A1(net3427),
    .S(_03252_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(net1797),
    .A1(net3558),
    .S(_03252_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _09264_ (.A0(net1922),
    .A1(net3496),
    .S(_03252_),
    .X(_00465_));
 sky130_fd_sc_hd__and2b_1 _09265_ (.A_N(net1545),
    .B(net1341),
    .X(_03253_));
 sky130_fd_sc_hd__and4bb_4 _09266_ (.A_N(net2407),
    .B_N(net1893),
    .C(net2787),
    .D(net1537),
    .X(_03254_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(net2664),
    .A1(net2368),
    .S(_03254_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _09268_ (.A0(net1705),
    .A1(net1875),
    .S(_03254_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(net1817),
    .A1(net2327),
    .S(_03254_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _09270_ (.A0(net1849),
    .A1(net1682),
    .S(_03254_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _09271_ (.A0(net2307),
    .A1(net2033),
    .S(_03254_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _09272_ (.A0(net2501),
    .A1(net2087),
    .S(_03254_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(net2536),
    .A1(net1797),
    .S(_03254_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _09274_ (.A0(net1361),
    .A1(net1922),
    .S(_03254_),
    .X(_00457_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(_03247_),
    .B(net2787),
    .Y(_03255_));
 sky130_fd_sc_hd__mux2_1 _09276_ (.A0(net2368),
    .A1(net1777),
    .S(net2788),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(net1875),
    .A1(net3037),
    .S(net2788),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _09278_ (.A0(net2327),
    .A1(net1801),
    .S(net2788),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(net1681),
    .A1(net1168),
    .S(net2788),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _09280_ (.A0(net2033),
    .A1(net1737),
    .S(net2788),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(net2087),
    .A1(net1786),
    .S(net2788),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _09282_ (.A0(net1797),
    .A1(net815),
    .S(net2788),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(net1921),
    .A1(net1118),
    .S(net2788),
    .X(_00449_));
 sky130_fd_sc_hd__nand2_8 _09284_ (.A(_03249_),
    .B(net2787),
    .Y(_03256_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(net2368),
    .A1(net1853),
    .S(_03256_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _09286_ (.A0(net1875),
    .A1(net2221),
    .S(_03256_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(net2327),
    .A1(net2114),
    .S(_03256_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(net1682),
    .A1(net3070),
    .S(_03256_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(net2033),
    .A1(net2231),
    .S(_03256_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _09290_ (.A0(net2087),
    .A1(net1733),
    .S(_03256_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(net1797),
    .A1(net1950),
    .S(_03256_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _09292_ (.A0(net1922),
    .A1(net2158),
    .S(_03256_),
    .X(_00441_));
 sky130_fd_sc_hd__nand2_4 _09293_ (.A(_03251_),
    .B(net2787),
    .Y(_03257_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(net2368),
    .A1(net752),
    .S(_03257_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(net1875),
    .A1(net2152),
    .S(_03257_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _09296_ (.A0(net2327),
    .A1(net2351),
    .S(_03257_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(net1682),
    .A1(net2345),
    .S(_03257_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(net2033),
    .A1(net2339),
    .S(_03257_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(net2087),
    .A1(net2068),
    .S(_03257_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _09300_ (.A0(net1797),
    .A1(net1241),
    .S(_03257_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(net1922),
    .A1(net1913),
    .S(_03257_),
    .X(_00433_));
 sky130_fd_sc_hd__and2_4 _09302_ (.A(net1341),
    .B(net1545),
    .X(_03258_));
 sky130_fd_sc_hd__nand2_1 _09303_ (.A(net1341),
    .B(net1545),
    .Y(_03259_));
 sky130_fd_sc_hd__and4bb_4 _09304_ (.A_N(net2407),
    .B_N(net1893),
    .C(_03258_),
    .D(net1537),
    .X(_03260_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(net2507),
    .A1(net2368),
    .S(_03260_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(net2415),
    .A1(net1875),
    .S(_03260_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(net1841),
    .A1(net2327),
    .S(_03260_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _09308_ (.A0(net2524),
    .A1(net1682),
    .S(_03260_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(net2530),
    .A1(net2033),
    .S(_03260_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(net1729),
    .A1(net2087),
    .S(_03260_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(net2542),
    .A1(net1797),
    .S(_03260_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(net2041),
    .A1(net1922),
    .S(_03260_),
    .X(_00425_));
 sky130_fd_sc_hd__nand2_4 _09313_ (.A(_03247_),
    .B(_03258_),
    .Y(_03261_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(net2367),
    .A1(net2686),
    .S(_03261_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(net1874),
    .A1(net1164),
    .S(_03261_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(net2326),
    .A1(net2678),
    .S(_03261_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(net1682),
    .A1(net3012),
    .S(_03261_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(net2032),
    .A1(net2972),
    .S(_03261_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(net2086),
    .A1(net2674),
    .S(_03261_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(net1796),
    .A1(net2682),
    .S(_03261_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(net1922),
    .A1(net2144),
    .S(_03261_),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_4 _09322_ (.A(_03249_),
    .B(_03258_),
    .Y(_03262_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(net2368),
    .A1(net3056),
    .S(_03262_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(net1875),
    .A1(net1917),
    .S(_03262_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(net2327),
    .A1(net2123),
    .S(_03262_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _09326_ (.A0(net1682),
    .A1(net2091),
    .S(_03262_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(net2033),
    .A1(net1833),
    .S(_03262_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _09328_ (.A0(net2087),
    .A1(net893),
    .S(_03262_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(net1797),
    .A1(net2106),
    .S(_03262_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(net1922),
    .A1(net3321),
    .S(_03262_),
    .X(_00409_));
 sky130_fd_sc_hd__and2_1 _09331_ (.A(net1198),
    .B(net1021),
    .X(_03263_));
 sky130_fd_sc_hd__a31o_1 _09332_ (.A1(net1580),
    .A2(net1198),
    .A3(net1021),
    .B1(net1245),
    .X(_00408_));
 sky130_fd_sc_hd__or3b_4 _09333_ (.A(net1580),
    .B(net1021),
    .C_N(net1596),
    .X(_03264_));
 sky130_fd_sc_hd__nor2_8 _09334_ (.A(_00666_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__a21o_1 _09335_ (.A1(net1537),
    .A2(_03264_),
    .B1(_03265_),
    .X(_00407_));
 sky130_fd_sc_hd__or3_1 _09336_ (.A(net360),
    .B(net1198),
    .C(net1022),
    .X(_03266_));
 sky130_fd_sc_hd__nor2_2 _09337_ (.A(_00667_),
    .B(net1023),
    .Y(_03267_));
 sky130_fd_sc_hd__a21o_1 _09338_ (.A1(net1337),
    .A2(net1023),
    .B1(net1024),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(net2368),
    .A1(net1065),
    .S(_03265_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _09340_ (.A0(net1875),
    .A1(net1059),
    .S(_03265_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _09341_ (.A0(net2327),
    .A1(net1029),
    .S(_03265_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(net1682),
    .A1(net1053),
    .S(_03265_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _09343_ (.A0(net2033),
    .A1(net1035),
    .S(_03265_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(net2087),
    .A1(net1041),
    .S(_03265_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(net1797),
    .A1(net1047),
    .S(_03265_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(net1922),
    .A1(net1071),
    .S(_03265_),
    .X(_00398_));
 sky130_fd_sc_hd__nand2_1 _09347_ (.A(_03243_),
    .B(_03265_),
    .Y(_03268_));
 sky130_fd_sc_hd__and3_1 _09348_ (.A(net1545),
    .B(_03243_),
    .C(_03265_),
    .X(_03269_));
 sky130_fd_sc_hd__o22a_1 _09349_ (.A1(_03259_),
    .A2(_03268_),
    .B1(net1546),
    .B2(net1341),
    .X(_00397_));
 sky130_fd_sc_hd__a21oi_1 _09350_ (.A1(_03243_),
    .A2(_03265_),
    .B1(net1545),
    .Y(_03270_));
 sky130_fd_sc_hd__nor2_1 _09351_ (.A(net1546),
    .B(net336),
    .Y(_00396_));
 sky130_fd_sc_hd__and2_1 _09352_ (.A(net1893),
    .B(_03265_),
    .X(_03271_));
 sky130_fd_sc_hd__o21a_1 _09353_ (.A1(net1599),
    .A2(net1894),
    .B1(_03268_),
    .X(_00395_));
 sky130_fd_sc_hd__nor2_1 _09354_ (.A(net1893),
    .B(_03265_),
    .Y(_03272_));
 sky130_fd_sc_hd__nor2_1 _09355_ (.A(net1894),
    .B(net455),
    .Y(_00394_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(net1377),
    .A1(net9),
    .S(net1024),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(net1389),
    .A1(net8),
    .S(net1024),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(net2287),
    .A1(net7),
    .S(net1024),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _09359_ (.A0(net1014),
    .A1(net6),
    .S(net1024),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(net1018),
    .A1(net5),
    .S(net1024),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(net1554),
    .A1(net4),
    .S(net1024),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(net1564),
    .A1(net3),
    .S(net1024),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _09363_ (.A0(net1373),
    .A1(net2),
    .S(net1024),
    .X(_00386_));
 sky130_fd_sc_hd__and3_1 _09364_ (.A(net1520),
    .B(net1444),
    .C(net1024),
    .X(_03273_));
 sky130_fd_sc_hd__a21oi_1 _09365_ (.A1(net1460),
    .A2(net1521),
    .B1(net1621),
    .Y(_03274_));
 sky130_fd_sc_hd__a21oi_1 _09366_ (.A1(net1622),
    .A2(net1521),
    .B1(net401),
    .Y(_00385_));
 sky130_fd_sc_hd__xor2_1 _09367_ (.A(net1460),
    .B(net1521),
    .X(_00384_));
 sky130_fd_sc_hd__a21oi_1 _09368_ (.A1(net1444),
    .A2(net1024),
    .B1(net1520),
    .Y(_03275_));
 sky130_fd_sc_hd__nor2_1 _09369_ (.A(net3368),
    .B(net389),
    .Y(_00383_));
 sky130_fd_sc_hd__xor2_1 _09370_ (.A(net1444),
    .B(net1024),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _09371_ (.A(net421),
    .B(net462),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_1 _09372_ (.A1(net971),
    .A2(net1898),
    .B1(net462),
    .B2(net421),
    .X(_03277_));
 sky130_fd_sc_hd__and3_1 _09373_ (.A(net971),
    .B(net1898),
    .C(net462),
    .X(_03278_));
 sky130_fd_sc_hd__a21bo_1 _09374_ (.A1(net421),
    .A2(_03278_),
    .B1_N(_03277_),
    .X(_03279_));
 sky130_fd_sc_hd__nand2_1 _09375_ (.A(net1381),
    .B(net1747),
    .Y(_03280_));
 sky130_fd_sc_hd__xor2_1 _09376_ (.A(_03279_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__and4_1 _09377_ (.A(net971),
    .B(net2225),
    .C(net1898),
    .D(net462),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_1 _09378_ (.A1(net2225),
    .A2(net1898),
    .B1(net462),
    .B2(net971),
    .X(_03283_));
 sky130_fd_sc_hd__inv_2 _09379_ (.A(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__and4b_1 _09380_ (.A_N(_03282_),
    .B(_03283_),
    .C(net421),
    .D(net1747),
    .X(_03285_));
 sky130_fd_sc_hd__o21ai_2 _09381_ (.A1(_03282_),
    .A2(_03285_),
    .B1(_03281_),
    .Y(_03286_));
 sky130_fd_sc_hd__or3_1 _09382_ (.A(_03281_),
    .B(_03282_),
    .C(_03285_),
    .X(_03287_));
 sky130_fd_sc_hd__nand2_1 _09383_ (.A(_03286_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__o2bb2a_1 _09384_ (.A1_N(net421),
    .A2_N(net1747),
    .B1(_03282_),
    .B2(_03284_),
    .X(_03289_));
 sky130_fd_sc_hd__or2_1 _09385_ (.A(_03285_),
    .B(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__nand4_1 _09386_ (.A(net2225),
    .B(net986),
    .C(net1898),
    .D(net462),
    .Y(_03291_));
 sky130_fd_sc_hd__a22o_1 _09387_ (.A1(net986),
    .A2(net1898),
    .B1(net462),
    .B2(net2225),
    .X(_03292_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(net971),
    .B(net1747),
    .Y(_03294_));
 sky130_fd_sc_hd__o21ai_1 _09390_ (.A1(_03293_),
    .A2(_03294_),
    .B1(_03291_),
    .Y(_03295_));
 sky130_fd_sc_hd__and2b_1 _09391_ (.A_N(_03290_),
    .B(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__and2b_1 _09392_ (.A_N(_03295_),
    .B(_03290_),
    .X(_03297_));
 sky130_fd_sc_hd__nor2_2 _09393_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_2 _09394_ (.A(net1381),
    .B(net722),
    .Y(_03299_));
 sky130_fd_sc_hd__a31oi_1 _09395_ (.A1(net1381),
    .A2(net722),
    .A3(_03298_),
    .B1(_03296_),
    .Y(_03300_));
 sky130_fd_sc_hd__or2_1 _09396_ (.A(_03288_),
    .B(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__nand2_1 _09397_ (.A(_03288_),
    .B(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__and2_1 _09398_ (.A(_03301_),
    .B(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_4 _09399_ (.A(_03298_),
    .B(_03299_),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_2 _09400_ (.A(_03293_),
    .B(_03294_),
    .Y(_03305_));
 sky130_fd_sc_hd__and4_1 _09401_ (.A(net986),
    .B(net827),
    .C(net1898),
    .D(net462),
    .X(_03306_));
 sky130_fd_sc_hd__a22oi_1 _09402_ (.A1(net827),
    .A2(net1898),
    .B1(net462),
    .B2(net986),
    .Y(_03307_));
 sky130_fd_sc_hd__or2_1 _09403_ (.A(_03306_),
    .B(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__nand2_1 _09404_ (.A(net2225),
    .B(net1747),
    .Y(_03309_));
 sky130_fd_sc_hd__o21ba_1 _09405_ (.A1(_03308_),
    .A2(_03309_),
    .B1_N(_03306_),
    .X(_03310_));
 sky130_fd_sc_hd__xnor2_2 _09406_ (.A(_03305_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__a22oi_2 _09407_ (.A1(net421),
    .A2(net722),
    .B1(net944),
    .B2(net1381),
    .Y(_03312_));
 sky130_fd_sc_hd__and4_2 _09408_ (.A(net1381),
    .B(net421),
    .C(net722),
    .D(net944),
    .X(_03313_));
 sky130_fd_sc_hd__nor2_1 _09409_ (.A(_03312_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__o32a_2 _09410_ (.A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .B1(_03310_),
    .B2(_03305_),
    .X(_03315_));
 sky130_fd_sc_hd__and2b_1 _09411_ (.A_N(_03315_),
    .B(_03304_),
    .X(_03316_));
 sky130_fd_sc_hd__xnor2_4 _09412_ (.A(_03304_),
    .B(_03315_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _09413_ (.A1(_03313_),
    .A2(_03317_),
    .B1(_03316_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2b_1 _09414_ (.A_N(_03318_),
    .B(_03303_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2b_1 _09415_ (.A_N(_03303_),
    .B(_03318_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _09416_ (.A(_03319_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_4 _09417_ (.A(_03313_),
    .B(_03317_),
    .Y(_03322_));
 sky130_fd_sc_hd__xnor2_2 _09418_ (.A(_03311_),
    .B(_03314_),
    .Y(_03323_));
 sky130_fd_sc_hd__xnor2_1 _09419_ (.A(_03308_),
    .B(_03309_),
    .Y(_03324_));
 sky130_fd_sc_hd__and4_1 _09420_ (.A(net827),
    .B(net773),
    .C(net1898),
    .D(net462),
    .X(_03325_));
 sky130_fd_sc_hd__a22o_1 _09421_ (.A1(net773),
    .A2(net1898),
    .B1(net462),
    .B2(net827),
    .X(_03326_));
 sky130_fd_sc_hd__nand2b_2 _09422_ (.A_N(_03325_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_2 _09423_ (.A(net986),
    .B(net1747),
    .Y(_03328_));
 sky130_fd_sc_hd__a31o_1 _09424_ (.A1(net986),
    .A2(net1747),
    .A3(_03326_),
    .B1(_03325_),
    .X(_03329_));
 sky130_fd_sc_hd__and2b_1 _09425_ (.A_N(_03324_),
    .B(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__xor2_1 _09426_ (.A(_03324_),
    .B(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__a22o_1 _09427_ (.A1(net971),
    .A2(net722),
    .B1(net944),
    .B2(net421),
    .X(_03332_));
 sky130_fd_sc_hd__and4_1 _09428_ (.A(net421),
    .B(net971),
    .C(net722),
    .D(net944),
    .X(_03333_));
 sky130_fd_sc_hd__nand4_1 _09429_ (.A(net421),
    .B(net971),
    .C(net722),
    .D(net944),
    .Y(_03334_));
 sky130_fd_sc_hd__a22oi_1 _09430_ (.A1(net1381),
    .A2(net2148),
    .B1(_03332_),
    .B2(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__and4_1 _09431_ (.A(net1381),
    .B(net2148),
    .C(_03332_),
    .D(_03334_),
    .X(_03336_));
 sky130_fd_sc_hd__or2_1 _09432_ (.A(_03335_),
    .B(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__nor2_1 _09433_ (.A(_03331_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__o21ai_4 _09434_ (.A1(_03330_),
    .A2(_03338_),
    .B1(_03323_),
    .Y(_03339_));
 sky130_fd_sc_hd__or3_2 _09435_ (.A(_03323_),
    .B(_03330_),
    .C(_03338_),
    .X(_03340_));
 sky130_fd_sc_hd__o211ai_4 _09436_ (.A1(_03333_),
    .A2(_03336_),
    .B1(_03339_),
    .C1(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_2 _09437_ (.A(_03339_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand2b_1 _09438_ (.A_N(_03322_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nor2_1 _09439_ (.A(_03321_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__and2_1 _09440_ (.A(_03321_),
    .B(_03343_),
    .X(_03345_));
 sky130_fd_sc_hd__or2_1 _09441_ (.A(_03344_),
    .B(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__a211o_1 _09442_ (.A1(_03339_),
    .A2(_03340_),
    .B1(_03333_),
    .C1(_03336_),
    .X(_03347_));
 sky130_fd_sc_hd__xor2_1 _09443_ (.A(_03331_),
    .B(_03337_),
    .X(_03348_));
 sky130_fd_sc_hd__xnor2_4 _09444_ (.A(_03327_),
    .B(_03328_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand4_2 _09445_ (.A(net773),
    .B(net1590),
    .C(net1898),
    .D(net462),
    .Y(_03350_));
 sky130_fd_sc_hd__a22o_1 _09446_ (.A1(net1590),
    .A2(net1898),
    .B1(net462),
    .B2(net773),
    .X(_03351_));
 sky130_fd_sc_hd__nand4_2 _09447_ (.A(net827),
    .B(net1747),
    .C(_03350_),
    .D(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand2_2 _09448_ (.A(_03350_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__and2b_1 _09449_ (.A_N(_03349_),
    .B(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__a22o_1 _09450_ (.A1(net2225),
    .A2(net722),
    .B1(net944),
    .B2(net971),
    .X(_03355_));
 sky130_fd_sc_hd__nand4_4 _09451_ (.A(net971),
    .B(net2225),
    .C(net722),
    .D(net944),
    .Y(_03356_));
 sky130_fd_sc_hd__nand4_4 _09452_ (.A(net421),
    .B(net2148),
    .C(_03355_),
    .D(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__a22o_1 _09453_ (.A1(net2950),
    .A2(net2148),
    .B1(_03355_),
    .B2(_03356_),
    .X(_03358_));
 sky130_fd_sc_hd__nand2_2 _09454_ (.A(_03357_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__xor2_4 _09455_ (.A(_03349_),
    .B(_03353_),
    .X(_03360_));
 sky130_fd_sc_hd__nor2_1 _09456_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__o21a_2 _09457_ (.A1(_03354_),
    .A2(_03361_),
    .B1(_03348_),
    .X(_03362_));
 sky130_fd_sc_hd__nor3_2 _09458_ (.A(_03348_),
    .B(_03354_),
    .C(_03361_),
    .Y(_03363_));
 sky130_fd_sc_hd__a211oi_4 _09459_ (.A1(_03356_),
    .A2(_03357_),
    .B1(_03362_),
    .C1(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__o211ai_4 _09460_ (.A1(_03362_),
    .A2(_03364_),
    .B1(_03341_),
    .C1(_03347_),
    .Y(_03365_));
 sky130_fd_sc_hd__xor2_4 _09461_ (.A(_03322_),
    .B(_03342_),
    .X(_03366_));
 sky130_fd_sc_hd__or2_1 _09462_ (.A(_03365_),
    .B(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__a211o_1 _09463_ (.A1(_03341_),
    .A2(_03347_),
    .B1(_03362_),
    .C1(_03364_),
    .X(_03368_));
 sky130_fd_sc_hd__nand2_1 _09464_ (.A(_03365_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__inv_2 _09465_ (.A(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o211ai_1 _09466_ (.A1(_03362_),
    .A2(_03363_),
    .B1(_03356_),
    .C1(_03357_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2b_1 _09467_ (.A_N(_03364_),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__xor2_4 _09468_ (.A(_03359_),
    .B(_03360_),
    .X(_03373_));
 sky130_fd_sc_hd__a22o_1 _09469_ (.A1(net827),
    .A2(net1747),
    .B1(_03350_),
    .B2(_03351_),
    .X(_03374_));
 sky130_fd_sc_hd__and4_1 _09470_ (.A(net773),
    .B(net1590),
    .C(net2027),
    .D(net1747),
    .X(_03375_));
 sky130_fd_sc_hd__nand3_1 _09471_ (.A(_03352_),
    .B(_03374_),
    .C(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__and4_1 _09472_ (.A(net2225),
    .B(net986),
    .C(net722),
    .D(net944),
    .X(_03377_));
 sky130_fd_sc_hd__a22o_1 _09473_ (.A1(net2517),
    .A2(net722),
    .B1(net944),
    .B2(net2225),
    .X(_03378_));
 sky130_fd_sc_hd__and2b_1 _09474_ (.A_N(_03377_),
    .B(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__nand2_1 _09475_ (.A(net971),
    .B(net2148),
    .Y(_03380_));
 sky130_fd_sc_hd__xnor2_2 _09476_ (.A(_03379_),
    .B(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__a21o_1 _09477_ (.A1(_03352_),
    .A2(_03374_),
    .B1(_03375_),
    .X(_03382_));
 sky130_fd_sc_hd__and3_1 _09478_ (.A(_03376_),
    .B(_03381_),
    .C(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__a21boi_4 _09479_ (.A1(_03381_),
    .A2(_03382_),
    .B1_N(_03376_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2b_1 _09480_ (.A_N(_03384_),
    .B(_03373_),
    .Y(_03385_));
 sky130_fd_sc_hd__a31o_1 _09481_ (.A1(net971),
    .A2(net2148),
    .A3(_03378_),
    .B1(_03377_),
    .X(_03386_));
 sky130_fd_sc_hd__and3_2 _09482_ (.A(net1381),
    .B(net1809),
    .C(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__a21oi_1 _09483_ (.A1(net1381),
    .A2(net1809),
    .B1(_03386_),
    .Y(_03388_));
 sky130_fd_sc_hd__or2_2 _09484_ (.A(_03387_),
    .B(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__xor2_4 _09485_ (.A(_03373_),
    .B(_03384_),
    .X(_03390_));
 sky130_fd_sc_hd__o21ai_2 _09486_ (.A1(_03389_),
    .A2(_03390_),
    .B1(_03385_),
    .Y(_03391_));
 sky130_fd_sc_hd__and2b_1 _09487_ (.A_N(_03372_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__xnor2_2 _09488_ (.A(_03372_),
    .B(_03391_),
    .Y(_03393_));
 sky130_fd_sc_hd__and2_1 _09489_ (.A(_03387_),
    .B(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__o21a_1 _09490_ (.A1(_03392_),
    .A2(_03394_),
    .B1(_03370_),
    .X(_03395_));
 sky130_fd_sc_hd__xnor2_4 _09491_ (.A(_03387_),
    .B(_03393_),
    .Y(_03396_));
 sky130_fd_sc_hd__xnor2_4 _09492_ (.A(_03389_),
    .B(_03390_),
    .Y(_03397_));
 sky130_fd_sc_hd__a21oi_1 _09493_ (.A1(_03376_),
    .A2(_03382_),
    .B1(_03381_),
    .Y(_03398_));
 sky130_fd_sc_hd__a22o_1 _09494_ (.A1(net827),
    .A2(net722),
    .B1(net944),
    .B2(net2517),
    .X(_03399_));
 sky130_fd_sc_hd__nand4_1 _09495_ (.A(net986),
    .B(net827),
    .C(net722),
    .D(net944),
    .Y(_03400_));
 sky130_fd_sc_hd__and2_1 _09496_ (.A(net2225),
    .B(net2148),
    .X(_03401_));
 sky130_fd_sc_hd__a21o_1 _09497_ (.A1(_03399_),
    .A2(_03400_),
    .B1(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__nand3_1 _09498_ (.A(_03399_),
    .B(_03400_),
    .C(_03401_),
    .Y(_03403_));
 sky130_fd_sc_hd__a22oi_1 _09499_ (.A1(net1590),
    .A2(net2027),
    .B1(net1747),
    .B2(net773),
    .Y(_03404_));
 sky130_fd_sc_hd__nor2_1 _09500_ (.A(_03375_),
    .B(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand3_1 _09501_ (.A(_03402_),
    .B(_03403_),
    .C(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__or3_1 _09502_ (.A(_03383_),
    .B(_03398_),
    .C(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__a21bo_1 _09503_ (.A1(_03399_),
    .A2(_03401_),
    .B1_N(_03400_),
    .X(_03408_));
 sky130_fd_sc_hd__and2_1 _09504_ (.A(net421),
    .B(net1809),
    .X(_03409_));
 sky130_fd_sc_hd__nor2_1 _09505_ (.A(_03408_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__and2_1 _09506_ (.A(_03408_),
    .B(_03409_),
    .X(_03411_));
 sky130_fd_sc_hd__nor2_1 _09507_ (.A(_03410_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(net1381),
    .B(net836),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _09509_ (.A(_03412_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__o21ai_1 _09510_ (.A1(_03383_),
    .A2(_03398_),
    .B1(_03406_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand3_1 _09511_ (.A(_03407_),
    .B(_03414_),
    .C(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_2 _09512_ (.A(_03407_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2b_1 _09513_ (.A_N(_03397_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__a31o_2 _09514_ (.A1(net1381),
    .A2(net836),
    .A3(_03412_),
    .B1(_03411_),
    .X(_03419_));
 sky130_fd_sc_hd__xnor2_4 _09515_ (.A(_03397_),
    .B(_03417_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21boi_4 _09516_ (.A1(_03419_),
    .A2(_03420_),
    .B1_N(_03418_),
    .Y(_03421_));
 sky130_fd_sc_hd__nor2_1 _09517_ (.A(_03396_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__xor2_4 _09518_ (.A(_03396_),
    .B(_03421_),
    .X(_03423_));
 sky130_fd_sc_hd__xnor2_2 _09519_ (.A(_03419_),
    .B(_03420_),
    .Y(_03424_));
 sky130_fd_sc_hd__a21o_1 _09520_ (.A1(_03407_),
    .A2(_03415_),
    .B1(_03414_),
    .X(_03425_));
 sky130_fd_sc_hd__a21o_1 _09521_ (.A1(_03402_),
    .A2(_03403_),
    .B1(_03405_),
    .X(_03426_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(net1590),
    .B(net1747),
    .Y(_03427_));
 sky130_fd_sc_hd__a22oi_1 _09523_ (.A1(net773),
    .A2(net722),
    .B1(net2394),
    .B2(net827),
    .Y(_03428_));
 sky130_fd_sc_hd__a22o_1 _09524_ (.A1(net773),
    .A2(net2389),
    .B1(net2394),
    .B2(net827),
    .X(_03429_));
 sky130_fd_sc_hd__and4_1 _09525_ (.A(net827),
    .B(net773),
    .C(net722),
    .D(net2394),
    .X(_03430_));
 sky130_fd_sc_hd__and4b_1 _09526_ (.A_N(_03430_),
    .B(net2148),
    .C(net986),
    .D(_03429_),
    .X(_03431_));
 sky130_fd_sc_hd__o2bb2a_1 _09527_ (.A1_N(net986),
    .A2_N(net2148),
    .B1(_03428_),
    .B2(_03430_),
    .X(_03432_));
 sky130_fd_sc_hd__nor3_1 _09528_ (.A(_03427_),
    .B(_03431_),
    .C(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand3_1 _09529_ (.A(_03406_),
    .B(_03426_),
    .C(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _09530_ (.A(net2950),
    .B(net2377),
    .Y(_03435_));
 sky130_fd_sc_hd__a31o_1 _09531_ (.A1(net986),
    .A2(net2148),
    .A3(_03429_),
    .B1(_03430_),
    .X(_03436_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(net971),
    .B(net1809),
    .Y(_03437_));
 sky130_fd_sc_hd__and3_1 _09533_ (.A(net971),
    .B(net1809),
    .C(_03436_),
    .X(_03438_));
 sky130_fd_sc_hd__xnor2_1 _09534_ (.A(_03436_),
    .B(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__and3_1 _09535_ (.A(net2950),
    .B(net836),
    .C(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__xnor2_1 _09536_ (.A(_03435_),
    .B(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__a21o_1 _09537_ (.A1(_03406_),
    .A2(_03426_),
    .B1(_03433_),
    .X(_03442_));
 sky130_fd_sc_hd__nand3_1 _09538_ (.A(_03434_),
    .B(_03441_),
    .C(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_1 _09539_ (.A(_03434_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand3_1 _09540_ (.A(_03416_),
    .B(_03425_),
    .C(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__a21o_1 _09541_ (.A1(_03416_),
    .A2(_03425_),
    .B1(_03444_),
    .X(_03446_));
 sky130_fd_sc_hd__o211ai_2 _09542_ (.A1(_03438_),
    .A2(_03440_),
    .B1(_03445_),
    .C1(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_03445_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__and2b_1 _09544_ (.A_N(_03424_),
    .B(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__xnor2_2 _09545_ (.A(_03424_),
    .B(_03448_),
    .Y(_03450_));
 sky130_fd_sc_hd__a211o_1 _09546_ (.A1(_03445_),
    .A2(_03446_),
    .B1(_03438_),
    .C1(_03440_),
    .X(_03451_));
 sky130_fd_sc_hd__a21o_1 _09547_ (.A1(_03434_),
    .A2(_03442_),
    .B1(_03441_),
    .X(_03452_));
 sky130_fd_sc_hd__nand2_1 _09548_ (.A(net971),
    .B(net836),
    .Y(_03453_));
 sky130_fd_sc_hd__and4_1 _09549_ (.A(net773),
    .B(net1590),
    .C(net2389),
    .D(net944),
    .X(_03454_));
 sky130_fd_sc_hd__nand2_1 _09550_ (.A(net827),
    .B(net2148),
    .Y(_03455_));
 sky130_fd_sc_hd__a22oi_2 _09551_ (.A1(net1590),
    .A2(net2389),
    .B1(net944),
    .B2(net773),
    .Y(_03456_));
 sky130_fd_sc_hd__nor2_1 _09552_ (.A(_03454_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__o21bai_1 _09553_ (.A1(_03455_),
    .A2(_03456_),
    .B1_N(_03454_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(net2225),
    .B(net1809),
    .Y(_03459_));
 sky130_fd_sc_hd__and3_1 _09555_ (.A(net2225),
    .B(net1809),
    .C(_03458_),
    .X(_03460_));
 sky130_fd_sc_hd__xnor2_1 _09556_ (.A(_03458_),
    .B(_03459_),
    .Y(_03461_));
 sky130_fd_sc_hd__xnor2_1 _09557_ (.A(_03453_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__o21a_1 _09558_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_03427_),
    .X(_03463_));
 sky130_fd_sc_hd__nor2_1 _09559_ (.A(_03433_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__and2_1 _09560_ (.A(_03462_),
    .B(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__and3_1 _09561_ (.A(_03443_),
    .B(_03452_),
    .C(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__a31o_1 _09562_ (.A1(net2511),
    .A2(net836),
    .A3(_03461_),
    .B1(_03460_),
    .X(_03467_));
 sky130_fd_sc_hd__inv_2 _09563_ (.A(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__a21oi_1 _09564_ (.A1(_03443_),
    .A2(_03452_),
    .B1(_03465_),
    .Y(_03469_));
 sky130_fd_sc_hd__nor3_1 _09565_ (.A(_03466_),
    .B(_03468_),
    .C(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__or3_1 _09566_ (.A(_03466_),
    .B(_03468_),
    .C(_03469_),
    .X(_03471_));
 sky130_fd_sc_hd__o211a_1 _09567_ (.A1(_03466_),
    .A2(_03470_),
    .B1(_03447_),
    .C1(_03451_),
    .X(_03472_));
 sky130_fd_sc_hd__a211o_1 _09568_ (.A1(_03447_),
    .A2(_03451_),
    .B1(_03466_),
    .C1(_03470_),
    .X(_03473_));
 sky130_fd_sc_hd__o21ai_1 _09569_ (.A1(_03466_),
    .A2(_03469_),
    .B1(_03468_),
    .Y(_03474_));
 sky130_fd_sc_hd__xnor2_1 _09570_ (.A(_03462_),
    .B(_03464_),
    .Y(_03475_));
 sky130_fd_sc_hd__xnor2_1 _09571_ (.A(_03455_),
    .B(_03457_),
    .Y(_03476_));
 sky130_fd_sc_hd__and4_1 _09572_ (.A(net1676),
    .B(net1590),
    .C(net944),
    .D(net2148),
    .X(_03477_));
 sky130_fd_sc_hd__inv_2 _09573_ (.A(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__a21oi_1 _09574_ (.A1(net986),
    .A2(net1809),
    .B1(_03477_),
    .Y(_03479_));
 sky130_fd_sc_hd__and3_1 _09575_ (.A(net986),
    .B(net1809),
    .C(_03477_),
    .X(_03480_));
 sky130_fd_sc_hd__nor2_1 _09576_ (.A(_03479_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(net2225),
    .B(net836),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor2_1 _09578_ (.A(_03481_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(_03476_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nor2_1 _09580_ (.A(_03475_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__a31o_1 _09581_ (.A1(net2225),
    .A2(net836),
    .A3(_03481_),
    .B1(_03480_),
    .X(_03486_));
 sky130_fd_sc_hd__xor2_1 _09582_ (.A(_03475_),
    .B(_03484_),
    .X(_03487_));
 sky130_fd_sc_hd__and2_1 _09583_ (.A(_03486_),
    .B(_03487_),
    .X(_03488_));
 sky130_fd_sc_hd__o211a_1 _09584_ (.A1(_03485_),
    .A2(_03488_),
    .B1(_03471_),
    .C1(_03474_),
    .X(_03489_));
 sky130_fd_sc_hd__a211o_1 _09585_ (.A1(_03471_),
    .A2(_03474_),
    .B1(_03485_),
    .C1(_03488_),
    .X(_03490_));
 sky130_fd_sc_hd__nand2b_1 _09586_ (.A_N(_03489_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__xnor2_1 _09587_ (.A(_03486_),
    .B(_03487_),
    .Y(_03492_));
 sky130_fd_sc_hd__xnor2_1 _09588_ (.A(_03476_),
    .B(_03483_),
    .Y(_03493_));
 sky130_fd_sc_hd__and4_1 _09589_ (.A(net986),
    .B(net827),
    .C(net1809),
    .D(net836),
    .X(_03494_));
 sky130_fd_sc_hd__inv_2 _09590_ (.A(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__a22o_1 _09591_ (.A1(net1590),
    .A2(net944),
    .B1(net2148),
    .B2(net773),
    .X(_03496_));
 sky130_fd_sc_hd__a22o_1 _09592_ (.A1(net827),
    .A2(net1809),
    .B1(net836),
    .B2(net986),
    .X(_03497_));
 sky130_fd_sc_hd__or4bb_1 _09593_ (.A(_03477_),
    .B(_03494_),
    .C_N(_03496_),
    .D_N(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__and2_1 _09594_ (.A(_03495_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__nor2_1 _09595_ (.A(_03493_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__xnor2_1 _09596_ (.A(_03493_),
    .B(_03499_),
    .Y(_03501_));
 sky130_fd_sc_hd__a22o_1 _09597_ (.A1(_03478_),
    .A2(_03496_),
    .B1(_03497_),
    .B2(_03495_),
    .X(_03502_));
 sky130_fd_sc_hd__and4_1 _09598_ (.A(net1699),
    .B(net1677),
    .C(net1809),
    .D(net836),
    .X(_03503_));
 sky130_fd_sc_hd__a22o_1 _09599_ (.A1(net1676),
    .A2(net1809),
    .B1(net836),
    .B2(net1698),
    .X(_03504_));
 sky130_fd_sc_hd__inv_2 _09600_ (.A(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__and4b_1 _09601_ (.A_N(_03503_),
    .B(_03504_),
    .C(net1590),
    .D(net2148),
    .X(_03506_));
 sky130_fd_sc_hd__or2_1 _09602_ (.A(_03503_),
    .B(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__and3_1 _09603_ (.A(_03498_),
    .B(_03502_),
    .C(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__o2bb2a_1 _09604_ (.A1_N(net1590),
    .A2_N(net2148),
    .B1(_03503_),
    .B2(_03505_),
    .X(_03509_));
 sky130_fd_sc_hd__nor2_1 _09605_ (.A(_03506_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__and4_1 _09606_ (.A(net1677),
    .B(net1590),
    .C(net1809),
    .D(net836),
    .X(_03511_));
 sky130_fd_sc_hd__and2_1 _09607_ (.A(_03510_),
    .B(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__a21oi_1 _09608_ (.A1(_03498_),
    .A2(_03502_),
    .B1(_03507_),
    .Y(_03513_));
 sky130_fd_sc_hd__nor2_1 _09609_ (.A(_03508_),
    .B(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__a21oi_1 _09610_ (.A1(_03512_),
    .A2(_03514_),
    .B1(_03508_),
    .Y(_03515_));
 sky130_fd_sc_hd__o21ba_1 _09611_ (.A1(_03501_),
    .A2(_03515_),
    .B1_N(_03500_),
    .X(_03516_));
 sky130_fd_sc_hd__nor2_2 _09612_ (.A(_03492_),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__a21o_1 _09613_ (.A1(_03490_),
    .A2(_03517_),
    .B1(_03489_),
    .X(_03518_));
 sky130_fd_sc_hd__a21o_1 _09614_ (.A1(_03473_),
    .A2(_03518_),
    .B1(_03472_),
    .X(_03519_));
 sky130_fd_sc_hd__a21o_2 _09615_ (.A1(_03450_),
    .A2(_03519_),
    .B1(_03449_),
    .X(_03520_));
 sky130_fd_sc_hd__a21oi_2 _09616_ (.A1(_03423_),
    .A2(_03520_),
    .B1(_03422_),
    .Y(_03521_));
 sky130_fd_sc_hd__nor3_1 _09617_ (.A(_03370_),
    .B(_03392_),
    .C(_03394_),
    .Y(_03522_));
 sky130_fd_sc_hd__or2_1 _09618_ (.A(_03395_),
    .B(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__o21ba_2 _09619_ (.A1(_03521_),
    .A2(_03523_),
    .B1_N(_03395_),
    .X(_03524_));
 sky130_fd_sc_hd__a211oi_4 _09620_ (.A1(_03365_),
    .A2(_03524_),
    .B1(_03366_),
    .C1(_03346_),
    .Y(_03525_));
 sky130_fd_sc_hd__o211a_1 _09621_ (.A1(_03366_),
    .A2(_03524_),
    .B1(_03367_),
    .C1(_03346_),
    .X(_03526_));
 sky130_fd_sc_hd__nor2_2 _09622_ (.A(_03525_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _09623_ (.A(net51),
    .B(net686),
    .Y(_03528_));
 sky130_fd_sc_hd__a22o_1 _09624_ (.A1(net830),
    .A2(net1991),
    .B1(net686),
    .B2(net51),
    .X(_03529_));
 sky130_fd_sc_hd__and3_1 _09625_ (.A(net830),
    .B(net1991),
    .C(net686),
    .X(_03530_));
 sky130_fd_sc_hd__a21bo_1 _09626_ (.A1(net51),
    .A2(_03530_),
    .B1_N(_03529_),
    .X(_03531_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(net1425),
    .B(net1845),
    .Y(_03532_));
 sky130_fd_sc_hd__xor2_1 _09628_ (.A(_03531_),
    .B(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__and4_1 _09629_ (.A(net830),
    .B(net2690),
    .C(net1991),
    .D(net686),
    .X(_03534_));
 sky130_fd_sc_hd__a22o_1 _09630_ (.A1(net1094),
    .A2(net1991),
    .B1(net686),
    .B2(net830),
    .X(_03535_));
 sky130_fd_sc_hd__inv_2 _09631_ (.A(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__and4b_1 _09632_ (.A_N(_03534_),
    .B(_03535_),
    .C(net51),
    .D(net1845),
    .X(_03537_));
 sky130_fd_sc_hd__o21ai_2 _09633_ (.A1(_03534_),
    .A2(_03537_),
    .B1(_03533_),
    .Y(_03538_));
 sky130_fd_sc_hd__or3_1 _09634_ (.A(_03533_),
    .B(_03534_),
    .C(_03537_),
    .X(_03539_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_03538_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o2bb2a_1 _09636_ (.A1_N(net51),
    .A2_N(net1845),
    .B1(_03534_),
    .B2(_03536_),
    .X(_03541_));
 sky130_fd_sc_hd__or2_1 _09637_ (.A(_03537_),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__nand4_1 _09638_ (.A(net1094),
    .B(net1172),
    .C(net1991),
    .D(net686),
    .Y(_03543_));
 sky130_fd_sc_hd__a22o_1 _09639_ (.A1(net1172),
    .A2(net1991),
    .B1(net686),
    .B2(net1094),
    .X(_03544_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(_03543_),
    .B(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(net830),
    .B(net1845),
    .Y(_03546_));
 sky130_fd_sc_hd__o21ai_1 _09642_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03543_),
    .Y(_03547_));
 sky130_fd_sc_hd__and2b_1 _09643_ (.A_N(_03542_),
    .B(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__and2b_1 _09644_ (.A_N(_03547_),
    .B(_03542_),
    .X(_03549_));
 sky130_fd_sc_hd__nor2_2 _09645_ (.A(_03548_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand2_2 _09646_ (.A(net1425),
    .B(net743),
    .Y(_03551_));
 sky130_fd_sc_hd__a31oi_1 _09647_ (.A1(net1425),
    .A2(net743),
    .A3(_03550_),
    .B1(_03548_),
    .Y(_03552_));
 sky130_fd_sc_hd__or2_1 _09648_ (.A(_03540_),
    .B(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__nand2_1 _09649_ (.A(_03540_),
    .B(_03552_),
    .Y(_03554_));
 sky130_fd_sc_hd__and2_1 _09650_ (.A(_03553_),
    .B(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__xnor2_4 _09651_ (.A(_03550_),
    .B(_03551_),
    .Y(_03556_));
 sky130_fd_sc_hd__xnor2_1 _09652_ (.A(_03545_),
    .B(_03546_),
    .Y(_03557_));
 sky130_fd_sc_hd__and4_1 _09653_ (.A(net1172),
    .B(net902),
    .C(net1991),
    .D(net2276),
    .X(_03558_));
 sky130_fd_sc_hd__a22oi_1 _09654_ (.A1(net902),
    .A2(net1991),
    .B1(net2276),
    .B2(net1172),
    .Y(_03559_));
 sky130_fd_sc_hd__or2_1 _09655_ (.A(_03558_),
    .B(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(net1094),
    .B(net1845),
    .Y(_03561_));
 sky130_fd_sc_hd__o21ba_1 _09657_ (.A1(_03560_),
    .A2(_03561_),
    .B1_N(_03558_),
    .X(_03562_));
 sky130_fd_sc_hd__xnor2_1 _09658_ (.A(_03557_),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__a22oi_2 _09659_ (.A1(net51),
    .A2(net743),
    .B1(net980),
    .B2(net1425),
    .Y(_03564_));
 sky130_fd_sc_hd__and4_2 _09660_ (.A(net1425),
    .B(net51),
    .C(net743),
    .D(net980),
    .X(_03565_));
 sky130_fd_sc_hd__nor2_1 _09661_ (.A(_03564_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__o32a_2 _09662_ (.A1(_03563_),
    .A2(_03564_),
    .A3(_03565_),
    .B1(_03562_),
    .B2(_03557_),
    .X(_03567_));
 sky130_fd_sc_hd__and2b_1 _09663_ (.A_N(_03567_),
    .B(_03556_),
    .X(_03568_));
 sky130_fd_sc_hd__xnor2_4 _09664_ (.A(_03556_),
    .B(_03567_),
    .Y(_03569_));
 sky130_fd_sc_hd__a21oi_1 _09665_ (.A1(_03565_),
    .A2(_03569_),
    .B1(_03568_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2b_2 _09666_ (.A_N(_03570_),
    .B(_03555_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand2b_1 _09667_ (.A_N(_03555_),
    .B(_03570_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(_03571_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__xnor2_4 _09669_ (.A(_03565_),
    .B(_03569_),
    .Y(_03574_));
 sky130_fd_sc_hd__xnor2_1 _09670_ (.A(_03563_),
    .B(_03566_),
    .Y(_03575_));
 sky130_fd_sc_hd__xnor2_1 _09671_ (.A(_03560_),
    .B(_03561_),
    .Y(_03576_));
 sky130_fd_sc_hd__and4_1 _09672_ (.A(net902),
    .B(net881),
    .C(net1991),
    .D(net686),
    .X(_03577_));
 sky130_fd_sc_hd__a22o_1 _09673_ (.A1(net881),
    .A2(net1991),
    .B1(net686),
    .B2(net902),
    .X(_03578_));
 sky130_fd_sc_hd__nand2b_1 _09674_ (.A_N(_03577_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _09675_ (.A(net1172),
    .B(net1845),
    .Y(_03580_));
 sky130_fd_sc_hd__a31o_1 _09676_ (.A1(net1172),
    .A2(net1845),
    .A3(_03578_),
    .B1(_03577_),
    .X(_03581_));
 sky130_fd_sc_hd__and2b_1 _09677_ (.A_N(_03576_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__xor2_1 _09678_ (.A(_03576_),
    .B(_03581_),
    .X(_03583_));
 sky130_fd_sc_hd__a22o_1 _09679_ (.A1(net830),
    .A2(net743),
    .B1(net980),
    .B2(net1345),
    .X(_03584_));
 sky130_fd_sc_hd__and4_1 _09680_ (.A(net51),
    .B(net830),
    .C(net743),
    .D(net980),
    .X(_03585_));
 sky130_fd_sc_hd__nand4_1 _09681_ (.A(net1345),
    .B(net830),
    .C(net2459),
    .D(net2464),
    .Y(_03586_));
 sky130_fd_sc_hd__a22oi_1 _09682_ (.A1(net1425),
    .A2(net2199),
    .B1(_03584_),
    .B2(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__and4_1 _09683_ (.A(net1425),
    .B(net2199),
    .C(_03584_),
    .D(_03586_),
    .X(_03588_));
 sky130_fd_sc_hd__or2_1 _09684_ (.A(_03587_),
    .B(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__nor2_1 _09685_ (.A(_03583_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__o21ai_2 _09686_ (.A1(_03582_),
    .A2(_03590_),
    .B1(_03575_),
    .Y(_03591_));
 sky130_fd_sc_hd__or3_2 _09687_ (.A(_03575_),
    .B(_03582_),
    .C(_03590_),
    .X(_03592_));
 sky130_fd_sc_hd__o211ai_4 _09688_ (.A1(_03585_),
    .A2(_03588_),
    .B1(_03591_),
    .C1(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_2 _09689_ (.A(_03591_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand2b_1 _09690_ (.A_N(_03574_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__nor2_1 _09691_ (.A(_03573_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__and2_1 _09692_ (.A(_03573_),
    .B(_03595_),
    .X(_03597_));
 sky130_fd_sc_hd__or2_1 _09693_ (.A(_03596_),
    .B(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__a211o_1 _09694_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03585_),
    .C1(_03588_),
    .X(_03599_));
 sky130_fd_sc_hd__xor2_1 _09695_ (.A(_03583_),
    .B(_03589_),
    .X(_03600_));
 sky130_fd_sc_hd__xnor2_2 _09696_ (.A(_03579_),
    .B(_03580_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand4_2 _09697_ (.A(net881),
    .B(net1607),
    .C(net1991),
    .D(net686),
    .Y(_03602_));
 sky130_fd_sc_hd__a22o_1 _09698_ (.A1(net1607),
    .A2(net1991),
    .B1(net686),
    .B2(net881),
    .X(_03603_));
 sky130_fd_sc_hd__nand4_2 _09699_ (.A(net902),
    .B(net1845),
    .C(_03602_),
    .D(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand2_1 _09700_ (.A(_03602_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__and2b_1 _09701_ (.A_N(_03601_),
    .B(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__a22o_1 _09702_ (.A1(net2690),
    .A2(net2459),
    .B1(net2464),
    .B2(net830),
    .X(_03607_));
 sky130_fd_sc_hd__nand4_4 _09703_ (.A(net3637),
    .B(net2690),
    .C(net2459),
    .D(net2464),
    .Y(_03608_));
 sky130_fd_sc_hd__nand4_2 _09704_ (.A(net51),
    .B(net2199),
    .C(_03607_),
    .D(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__a22o_1 _09705_ (.A1(net51),
    .A2(net2199),
    .B1(_03607_),
    .B2(_03608_),
    .X(_03610_));
 sky130_fd_sc_hd__nand2_1 _09706_ (.A(_03609_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__xor2_2 _09707_ (.A(_03601_),
    .B(_03605_),
    .X(_03612_));
 sky130_fd_sc_hd__nor2_1 _09708_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__o21a_2 _09709_ (.A1(_03606_),
    .A2(_03613_),
    .B1(_03600_),
    .X(_03614_));
 sky130_fd_sc_hd__nor3_1 _09710_ (.A(_03600_),
    .B(_03606_),
    .C(_03613_),
    .Y(_03615_));
 sky130_fd_sc_hd__a211oi_2 _09711_ (.A1(_03608_),
    .A2(_03609_),
    .B1(_03614_),
    .C1(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__o211ai_4 _09712_ (.A1(_03614_),
    .A2(_03616_),
    .B1(_03593_),
    .C1(_03599_),
    .Y(_03617_));
 sky130_fd_sc_hd__xor2_4 _09713_ (.A(_03574_),
    .B(_03594_),
    .X(_03618_));
 sky130_fd_sc_hd__or2_1 _09714_ (.A(_03617_),
    .B(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__a211o_1 _09715_ (.A1(_03593_),
    .A2(_03599_),
    .B1(_03614_),
    .C1(_03616_),
    .X(_03620_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_03617_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__inv_2 _09717_ (.A(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__o211ai_1 _09718_ (.A1(_03614_),
    .A2(_03615_),
    .B1(_03608_),
    .C1(_03609_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2b_1 _09719_ (.A_N(_03616_),
    .B(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__xor2_2 _09720_ (.A(_03611_),
    .B(_03612_),
    .X(_03625_));
 sky130_fd_sc_hd__a22o_1 _09721_ (.A1(net902),
    .A2(net1845),
    .B1(_03602_),
    .B2(_03603_),
    .X(_03626_));
 sky130_fd_sc_hd__and4_1 _09722_ (.A(net881),
    .B(net1607),
    .C(net686),
    .D(net1845),
    .X(_03627_));
 sky130_fd_sc_hd__nand3_1 _09723_ (.A(_03604_),
    .B(_03626_),
    .C(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__and4_1 _09724_ (.A(net1094),
    .B(net2846),
    .C(net743),
    .D(net980),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _09725_ (.A1(net2846),
    .A2(net743),
    .B1(net980),
    .B2(net1094),
    .X(_03630_));
 sky130_fd_sc_hd__and2b_1 _09726_ (.A_N(_03629_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nand2_1 _09727_ (.A(net830),
    .B(net2199),
    .Y(_03632_));
 sky130_fd_sc_hd__xnor2_1 _09728_ (.A(_03631_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__a21o_1 _09729_ (.A1(_03604_),
    .A2(_03626_),
    .B1(_03627_),
    .X(_03634_));
 sky130_fd_sc_hd__and3_1 _09730_ (.A(_03628_),
    .B(_03633_),
    .C(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__a21boi_1 _09731_ (.A1(_03633_),
    .A2(_03634_),
    .B1_N(_03628_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2b_1 _09732_ (.A_N(_03636_),
    .B(_03625_),
    .Y(_03637_));
 sky130_fd_sc_hd__a31o_1 _09733_ (.A1(net830),
    .A2(net2199),
    .A3(_03630_),
    .B1(_03629_),
    .X(_03638_));
 sky130_fd_sc_hd__and3_1 _09734_ (.A(net1425),
    .B(net1805),
    .C(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a21oi_1 _09735_ (.A1(net1425),
    .A2(net1805),
    .B1(_03638_),
    .Y(_03640_));
 sky130_fd_sc_hd__or2_2 _09736_ (.A(_03639_),
    .B(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__and2b_1 _09737_ (.A_N(_03625_),
    .B(_03636_),
    .X(_03642_));
 sky130_fd_sc_hd__xnor2_1 _09738_ (.A(_03625_),
    .B(_03636_),
    .Y(_03643_));
 sky130_fd_sc_hd__o21ai_2 _09739_ (.A1(_03641_),
    .A2(_03642_),
    .B1(_03637_),
    .Y(_03644_));
 sky130_fd_sc_hd__and2b_1 _09740_ (.A_N(_03624_),
    .B(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__xnor2_2 _09741_ (.A(_03624_),
    .B(_03644_),
    .Y(_03646_));
 sky130_fd_sc_hd__and2_1 _09742_ (.A(_03639_),
    .B(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__o21a_1 _09743_ (.A1(_03645_),
    .A2(_03647_),
    .B1(_03622_),
    .X(_03648_));
 sky130_fd_sc_hd__xnor2_2 _09744_ (.A(_03639_),
    .B(_03646_),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_2 _09745_ (.A(_03641_),
    .B(_03643_),
    .Y(_03650_));
 sky130_fd_sc_hd__a21oi_1 _09746_ (.A1(_03628_),
    .A2(_03634_),
    .B1(_03633_),
    .Y(_03651_));
 sky130_fd_sc_hd__a22o_1 _09747_ (.A1(net902),
    .A2(net743),
    .B1(net980),
    .B2(net1172),
    .X(_03652_));
 sky130_fd_sc_hd__nand4_2 _09748_ (.A(net1172),
    .B(net902),
    .C(net743),
    .D(net980),
    .Y(_03653_));
 sky130_fd_sc_hd__and2_1 _09749_ (.A(net2690),
    .B(net2199),
    .X(_03654_));
 sky130_fd_sc_hd__a21o_1 _09750_ (.A1(_03652_),
    .A2(_03653_),
    .B1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__nand3_1 _09751_ (.A(_03652_),
    .B(_03653_),
    .C(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__a22oi_1 _09752_ (.A1(net1607),
    .A2(net686),
    .B1(net1845),
    .B2(net881),
    .Y(_03657_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(_03627_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand3_2 _09754_ (.A(_03655_),
    .B(_03656_),
    .C(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__or3_1 _09755_ (.A(_03635_),
    .B(_03651_),
    .C(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__a21bo_1 _09756_ (.A1(_03652_),
    .A2(_03654_),
    .B1_N(_03653_),
    .X(_03661_));
 sky130_fd_sc_hd__and2_1 _09757_ (.A(net51),
    .B(net1805),
    .X(_03662_));
 sky130_fd_sc_hd__nor2_1 _09758_ (.A(_03661_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__and2_1 _09759_ (.A(_03661_),
    .B(_03662_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(_03663_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _09761_ (.A(net1425),
    .B(net2078),
    .Y(_03666_));
 sky130_fd_sc_hd__xnor2_1 _09762_ (.A(_03665_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__o21ai_2 _09763_ (.A1(_03635_),
    .A2(_03651_),
    .B1(_03659_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand3_1 _09764_ (.A(_03660_),
    .B(_03667_),
    .C(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _09765_ (.A(_03660_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_03650_),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__o21ba_1 _09767_ (.A1(_03663_),
    .A2(_03666_),
    .B1_N(_03664_),
    .X(_03672_));
 sky130_fd_sc_hd__xnor2_2 _09768_ (.A(_03650_),
    .B(_03670_),
    .Y(_03673_));
 sky130_fd_sc_hd__o21a_1 _09769_ (.A1(_03672_),
    .A2(_03673_),
    .B1(_03671_),
    .X(_03674_));
 sky130_fd_sc_hd__nor2_1 _09770_ (.A(_03649_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _09771_ (.A(_03649_),
    .B(_03674_),
    .Y(_03676_));
 sky130_fd_sc_hd__xnor2_2 _09772_ (.A(_03649_),
    .B(_03674_),
    .Y(_03677_));
 sky130_fd_sc_hd__xnor2_2 _09773_ (.A(_03672_),
    .B(_03673_),
    .Y(_03678_));
 sky130_fd_sc_hd__a21o_1 _09774_ (.A1(_03660_),
    .A2(_03668_),
    .B1(_03667_),
    .X(_03679_));
 sky130_fd_sc_hd__a21o_1 _09775_ (.A1(_03655_),
    .A2(_03656_),
    .B1(_03658_),
    .X(_03680_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(net1607),
    .B(net1845),
    .Y(_03681_));
 sky130_fd_sc_hd__a22oi_1 _09777_ (.A1(net881),
    .A2(net743),
    .B1(net980),
    .B2(net3430),
    .Y(_03682_));
 sky130_fd_sc_hd__a22o_1 _09778_ (.A1(net1751),
    .A2(net743),
    .B1(net980),
    .B2(net902),
    .X(_03683_));
 sky130_fd_sc_hd__and4_1 _09779_ (.A(net902),
    .B(net1751),
    .C(net743),
    .D(net980),
    .X(_03684_));
 sky130_fd_sc_hd__and4b_1 _09780_ (.A_N(_03684_),
    .B(net2199),
    .C(net1172),
    .D(_03683_),
    .X(_03685_));
 sky130_fd_sc_hd__o2bb2a_1 _09781_ (.A1_N(net1172),
    .A2_N(net2199),
    .B1(_03682_),
    .B2(_03684_),
    .X(_03686_));
 sky130_fd_sc_hd__nor3_1 _09782_ (.A(_03681_),
    .B(_03685_),
    .C(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand3_1 _09783_ (.A(_03659_),
    .B(_03680_),
    .C(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__nand2_1 _09784_ (.A(net51),
    .B(net2078),
    .Y(_03689_));
 sky130_fd_sc_hd__a31o_1 _09785_ (.A1(net1172),
    .A2(net2199),
    .A3(_03683_),
    .B1(_03684_),
    .X(_03690_));
 sky130_fd_sc_hd__nand2_1 _09786_ (.A(net830),
    .B(net1805),
    .Y(_03691_));
 sky130_fd_sc_hd__and3_1 _09787_ (.A(net830),
    .B(net1805),
    .C(_03690_),
    .X(_03692_));
 sky130_fd_sc_hd__xnor2_1 _09788_ (.A(_03690_),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__and3_1 _09789_ (.A(net51),
    .B(net2078),
    .C(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__xnor2_1 _09790_ (.A(_03689_),
    .B(_03693_),
    .Y(_03695_));
 sky130_fd_sc_hd__a21o_1 _09791_ (.A1(_03659_),
    .A2(_03680_),
    .B1(_03687_),
    .X(_03696_));
 sky130_fd_sc_hd__nand3_1 _09792_ (.A(_03688_),
    .B(_03695_),
    .C(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_1 _09793_ (.A(_03688_),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand3_1 _09794_ (.A(_03669_),
    .B(_03679_),
    .C(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21o_1 _09795_ (.A1(_03669_),
    .A2(_03679_),
    .B1(_03698_),
    .X(_03700_));
 sky130_fd_sc_hd__o211ai_2 _09796_ (.A1(_03692_),
    .A2(_03694_),
    .B1(_03699_),
    .C1(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__nand2_1 _09797_ (.A(_03699_),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__and2b_1 _09798_ (.A_N(_03678_),
    .B(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__xnor2_2 _09799_ (.A(_03678_),
    .B(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__a211o_1 _09800_ (.A1(_03699_),
    .A2(_03700_),
    .B1(_03692_),
    .C1(_03694_),
    .X(_03705_));
 sky130_fd_sc_hd__a21o_1 _09801_ (.A1(_03688_),
    .A2(_03696_),
    .B1(_03695_),
    .X(_03706_));
 sky130_fd_sc_hd__nand2_1 _09802_ (.A(net830),
    .B(net2078),
    .Y(_03707_));
 sky130_fd_sc_hd__and4_1 _09803_ (.A(net881),
    .B(net1607),
    .C(net743),
    .D(net980),
    .X(_03708_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(net902),
    .B(net2199),
    .Y(_03709_));
 sky130_fd_sc_hd__a22oi_2 _09805_ (.A1(net1607),
    .A2(net743),
    .B1(net980),
    .B2(net881),
    .Y(_03710_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_03708_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__o21bai_1 _09807_ (.A1(_03709_),
    .A2(_03710_),
    .B1_N(_03708_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _09808_ (.A(net2690),
    .B(net1805),
    .Y(_03713_));
 sky130_fd_sc_hd__and3_1 _09809_ (.A(net2690),
    .B(net1805),
    .C(_03712_),
    .X(_03714_));
 sky130_fd_sc_hd__xnor2_1 _09810_ (.A(_03712_),
    .B(_03713_),
    .Y(_03715_));
 sky130_fd_sc_hd__xnor2_1 _09811_ (.A(_03707_),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__o21a_1 _09812_ (.A1(_03685_),
    .A2(_03686_),
    .B1(_03681_),
    .X(_03717_));
 sky130_fd_sc_hd__nor2_1 _09813_ (.A(_03687_),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__and2_1 _09814_ (.A(_03716_),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__and3_1 _09815_ (.A(_03697_),
    .B(_03706_),
    .C(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__a31oi_2 _09816_ (.A1(net830),
    .A2(net2078),
    .A3(_03715_),
    .B1(_03714_),
    .Y(_03721_));
 sky130_fd_sc_hd__a21oi_1 _09817_ (.A1(_03697_),
    .A2(_03706_),
    .B1(_03719_),
    .Y(_03722_));
 sky130_fd_sc_hd__nor3_1 _09818_ (.A(_03720_),
    .B(_03721_),
    .C(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__or3_1 _09819_ (.A(_03720_),
    .B(_03721_),
    .C(_03722_),
    .X(_03724_));
 sky130_fd_sc_hd__o211a_1 _09820_ (.A1(_03720_),
    .A2(_03723_),
    .B1(_03701_),
    .C1(_03705_),
    .X(_03725_));
 sky130_fd_sc_hd__a211o_1 _09821_ (.A1(_03701_),
    .A2(_03705_),
    .B1(_03720_),
    .C1(_03723_),
    .X(_03726_));
 sky130_fd_sc_hd__o21ai_1 _09822_ (.A1(_03720_),
    .A2(_03722_),
    .B1(_03721_),
    .Y(_03727_));
 sky130_fd_sc_hd__xnor2_1 _09823_ (.A(_03716_),
    .B(_03718_),
    .Y(_03728_));
 sky130_fd_sc_hd__xnor2_1 _09824_ (.A(_03709_),
    .B(_03711_),
    .Y(_03729_));
 sky130_fd_sc_hd__and4_1 _09825_ (.A(net881),
    .B(net1607),
    .C(net980),
    .D(net2199),
    .X(_03730_));
 sky130_fd_sc_hd__inv_2 _09826_ (.A(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__a21oi_1 _09827_ (.A1(net1172),
    .A2(net1805),
    .B1(_03730_),
    .Y(_03732_));
 sky130_fd_sc_hd__and3_1 _09828_ (.A(net1172),
    .B(net1805),
    .C(_03730_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_1 _09829_ (.A(_03732_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(net2690),
    .B(net2078),
    .Y(_03735_));
 sky130_fd_sc_hd__xnor2_1 _09831_ (.A(_03734_),
    .B(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(_03729_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__nor2_1 _09833_ (.A(_03728_),
    .B(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__a31o_1 _09834_ (.A1(net2690),
    .A2(net2078),
    .A3(_03734_),
    .B1(_03733_),
    .X(_03739_));
 sky130_fd_sc_hd__xor2_1 _09835_ (.A(_03728_),
    .B(_03737_),
    .X(_03740_));
 sky130_fd_sc_hd__and2_1 _09836_ (.A(_03739_),
    .B(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__o211a_1 _09837_ (.A1(_03738_),
    .A2(_03741_),
    .B1(_03724_),
    .C1(_03727_),
    .X(_03742_));
 sky130_fd_sc_hd__a211o_1 _09838_ (.A1(_03724_),
    .A2(_03727_),
    .B1(_03738_),
    .C1(_03741_),
    .X(_03743_));
 sky130_fd_sc_hd__nand2b_1 _09839_ (.A_N(_03742_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__xnor2_1 _09840_ (.A(_03739_),
    .B(_03740_),
    .Y(_03745_));
 sky130_fd_sc_hd__xnor2_1 _09841_ (.A(_03729_),
    .B(_03736_),
    .Y(_03746_));
 sky130_fd_sc_hd__and4_1 _09842_ (.A(net1172),
    .B(net902),
    .C(net1805),
    .D(net2078),
    .X(_03747_));
 sky130_fd_sc_hd__inv_2 _09843_ (.A(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__a22o_1 _09844_ (.A1(net1607),
    .A2(net980),
    .B1(net2199),
    .B2(net881),
    .X(_03749_));
 sky130_fd_sc_hd__a22o_1 _09845_ (.A1(net902),
    .A2(net1805),
    .B1(net2078),
    .B2(net1172),
    .X(_03750_));
 sky130_fd_sc_hd__or4bb_1 _09846_ (.A(_03730_),
    .B(_03747_),
    .C_N(_03749_),
    .D_N(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(_03748_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand2b_1 _09848_ (.A_N(_03746_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__xor2_1 _09849_ (.A(_03746_),
    .B(_03752_),
    .X(_03754_));
 sky130_fd_sc_hd__a22o_1 _09850_ (.A1(_03731_),
    .A2(_03749_),
    .B1(_03750_),
    .B2(_03748_),
    .X(_03755_));
 sky130_fd_sc_hd__and4_1 _09851_ (.A(net1782),
    .B(net1752),
    .C(net1805),
    .D(net2078),
    .X(_03756_));
 sky130_fd_sc_hd__a22o_1 _09852_ (.A1(net1752),
    .A2(net1805),
    .B1(net2078),
    .B2(net1782),
    .X(_03757_));
 sky130_fd_sc_hd__inv_2 _09853_ (.A(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__and4b_1 _09854_ (.A_N(_03756_),
    .B(_03757_),
    .C(net1607),
    .D(net2199),
    .X(_03759_));
 sky130_fd_sc_hd__or2_1 _09855_ (.A(_03756_),
    .B(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__and3_1 _09856_ (.A(_03751_),
    .B(_03755_),
    .C(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__o2bb2a_1 _09857_ (.A1_N(net1607),
    .A2_N(net2199),
    .B1(_03756_),
    .B2(_03758_),
    .X(_03762_));
 sky130_fd_sc_hd__nor2_1 _09858_ (.A(_03759_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__and4_1 _09859_ (.A(net1752),
    .B(net1607),
    .C(net1805),
    .D(net2078),
    .X(_03764_));
 sky130_fd_sc_hd__and2_1 _09860_ (.A(_03763_),
    .B(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a21oi_1 _09861_ (.A1(_03751_),
    .A2(_03755_),
    .B1(_03760_),
    .Y(_03766_));
 sky130_fd_sc_hd__nor2_1 _09862_ (.A(_03761_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__a21oi_1 _09863_ (.A1(_03765_),
    .A2(_03767_),
    .B1(_03761_),
    .Y(_03768_));
 sky130_fd_sc_hd__or2_1 _09864_ (.A(_03754_),
    .B(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__a21oi_2 _09865_ (.A1(_03753_),
    .A2(_03769_),
    .B1(_03745_),
    .Y(_03770_));
 sky130_fd_sc_hd__a21o_1 _09866_ (.A1(_03743_),
    .A2(_03770_),
    .B1(_03742_),
    .X(_03771_));
 sky130_fd_sc_hd__a21o_1 _09867_ (.A1(_03726_),
    .A2(_03771_),
    .B1(_03725_),
    .X(_03772_));
 sky130_fd_sc_hd__a21o_1 _09868_ (.A1(_03704_),
    .A2(_03772_),
    .B1(_03703_),
    .X(_03773_));
 sky130_fd_sc_hd__a21o_1 _09869_ (.A1(_03676_),
    .A2(_03773_),
    .B1(_03675_),
    .X(_03774_));
 sky130_fd_sc_hd__or3_2 _09870_ (.A(_03622_),
    .B(_03645_),
    .C(_03647_),
    .X(_03775_));
 sky130_fd_sc_hd__nand2b_1 _09871_ (.A_N(_03648_),
    .B(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__a21oi_4 _09872_ (.A1(_03774_),
    .A2(_03775_),
    .B1(_03648_),
    .Y(_03777_));
 sky130_fd_sc_hd__a211oi_4 _09873_ (.A1(_03617_),
    .A2(_03777_),
    .B1(_03618_),
    .C1(_03598_),
    .Y(_03778_));
 sky130_fd_sc_hd__o211a_1 _09874_ (.A1(_03618_),
    .A2(_03777_),
    .B1(_03619_),
    .C1(_03598_),
    .X(_03779_));
 sky130_fd_sc_hd__nor2_2 _09875_ (.A(_03778_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(_03527_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_1 _09877_ (.A(net440),
    .B(net675),
    .Y(_03782_));
 sky130_fd_sc_hd__a22o_1 _09878_ (.A1(net932),
    .A2(net1857),
    .B1(net675),
    .B2(net440),
    .X(_03783_));
 sky130_fd_sc_hd__and3_1 _09879_ (.A(net440),
    .B(net1857),
    .C(net675),
    .X(_03784_));
 sky130_fd_sc_hd__a21bo_1 _09880_ (.A1(net932),
    .A2(_03784_),
    .B1_N(_03783_),
    .X(_03785_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(net1393),
    .B(net1870),
    .Y(_03786_));
 sky130_fd_sc_hd__xnor2_1 _09882_ (.A(_03785_),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__and4_1 _09883_ (.A(net932),
    .B(net2262),
    .C(net1857),
    .D(net675),
    .X(_03788_));
 sky130_fd_sc_hd__a22o_1 _09884_ (.A1(net2262),
    .A2(net1857),
    .B1(net675),
    .B2(net932),
    .X(_03789_));
 sky130_fd_sc_hd__inv_2 _09885_ (.A(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__and4b_1 _09886_ (.A_N(_03788_),
    .B(_03789_),
    .C(net440),
    .D(net1870),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_1 _09887_ (.A(_03788_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__or2_1 _09888_ (.A(_03787_),
    .B(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(_03787_),
    .B(_03792_),
    .Y(_03794_));
 sky130_fd_sc_hd__o2bb2a_1 _09890_ (.A1_N(net440),
    .A2_N(net1870),
    .B1(_03788_),
    .B2(_03790_),
    .X(_03795_));
 sky130_fd_sc_hd__or2_1 _09891_ (.A(_03791_),
    .B(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__nand4_1 _09892_ (.A(net2262),
    .B(net1879),
    .C(net1857),
    .D(net675),
    .Y(_03797_));
 sky130_fd_sc_hd__a22o_1 _09893_ (.A1(net1879),
    .A2(net1857),
    .B1(net675),
    .B2(net2262),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_1 _09894_ (.A(_03797_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__nand2_1 _09895_ (.A(net932),
    .B(net1870),
    .Y(_03800_));
 sky130_fd_sc_hd__o21ai_1 _09896_ (.A1(_03799_),
    .A2(_03800_),
    .B1(_03797_),
    .Y(_03801_));
 sky130_fd_sc_hd__and2b_1 _09897_ (.A_N(_03796_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__and2b_1 _09898_ (.A_N(_03801_),
    .B(_03796_),
    .X(_03803_));
 sky130_fd_sc_hd__nor2_1 _09899_ (.A(_03802_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(net1393),
    .B(net746),
    .Y(_03805_));
 sky130_fd_sc_hd__a31oi_2 _09901_ (.A1(net1393),
    .A2(net746),
    .A3(_03804_),
    .B1(_03802_),
    .Y(_03806_));
 sky130_fd_sc_hd__or2_1 _09902_ (.A(_03794_),
    .B(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2_1 _09903_ (.A(_03794_),
    .B(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__and2_1 _09904_ (.A(_03807_),
    .B(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__xnor2_1 _09905_ (.A(_03804_),
    .B(_03805_),
    .Y(_03810_));
 sky130_fd_sc_hd__xnor2_1 _09906_ (.A(_03799_),
    .B(_03800_),
    .Y(_03811_));
 sky130_fd_sc_hd__and4_1 _09907_ (.A(net1879),
    .B(net863),
    .C(net1857),
    .D(net675),
    .X(_03812_));
 sky130_fd_sc_hd__a22o_1 _09908_ (.A1(net863),
    .A2(net1857),
    .B1(net675),
    .B2(net1879),
    .X(_03813_));
 sky130_fd_sc_hd__nand2b_1 _09909_ (.A_N(_03812_),
    .B(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand2_1 _09910_ (.A(net2262),
    .B(net1870),
    .Y(_03815_));
 sky130_fd_sc_hd__a31o_1 _09911_ (.A1(net2262),
    .A2(net1870),
    .A3(_03813_),
    .B1(_03812_),
    .X(_03816_));
 sky130_fd_sc_hd__nand2b_1 _09912_ (.A_N(_03811_),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__xor2_1 _09913_ (.A(_03811_),
    .B(_03816_),
    .X(_03818_));
 sky130_fd_sc_hd__a22oi_1 _09914_ (.A1(net440),
    .A2(net746),
    .B1(net875),
    .B2(net1393),
    .Y(_03819_));
 sky130_fd_sc_hd__and4_1 _09915_ (.A(net1393),
    .B(net440),
    .C(net746),
    .D(net875),
    .X(_03820_));
 sky130_fd_sc_hd__nor2_1 _09916_ (.A(_03819_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__o31a_1 _09917_ (.A1(_03818_),
    .A2(_03819_),
    .A3(_03820_),
    .B1(_03817_),
    .X(_03822_));
 sky130_fd_sc_hd__and2b_1 _09918_ (.A_N(_03822_),
    .B(_03810_),
    .X(_03823_));
 sky130_fd_sc_hd__xnor2_1 _09919_ (.A(_03810_),
    .B(_03822_),
    .Y(_03824_));
 sky130_fd_sc_hd__a21oi_1 _09920_ (.A1(_03820_),
    .A2(_03824_),
    .B1(_03823_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2b_1 _09921_ (.A_N(_03825_),
    .B(_03809_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2b_1 _09922_ (.A_N(_03809_),
    .B(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _09923_ (.A(_03826_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _09924_ (.A(_03820_),
    .B(_03824_),
    .Y(_03829_));
 sky130_fd_sc_hd__xnor2_1 _09925_ (.A(_03818_),
    .B(_03821_),
    .Y(_03830_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_03814_),
    .B(_03815_),
    .Y(_03831_));
 sky130_fd_sc_hd__and4_1 _09927_ (.A(net863),
    .B(net812),
    .C(net1857),
    .D(net2798),
    .X(_03832_));
 sky130_fd_sc_hd__a22o_1 _09928_ (.A1(net812),
    .A2(net1857),
    .B1(net2798),
    .B2(net863),
    .X(_03833_));
 sky130_fd_sc_hd__nand2b_1 _09929_ (.A_N(_03832_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(net1879),
    .B(net1870),
    .Y(_03835_));
 sky130_fd_sc_hd__a31o_1 _09931_ (.A1(net1879),
    .A2(net1870),
    .A3(_03833_),
    .B1(_03832_),
    .X(_03836_));
 sky130_fd_sc_hd__and2b_1 _09932_ (.A_N(_03831_),
    .B(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__xor2_1 _09933_ (.A(_03831_),
    .B(_03836_),
    .X(_03838_));
 sky130_fd_sc_hd__a22o_1 _09934_ (.A1(net932),
    .A2(net2869),
    .B1(net875),
    .B2(net440),
    .X(_03839_));
 sky130_fd_sc_hd__and4_1 _09935_ (.A(net3682),
    .B(net932),
    .C(net2869),
    .D(net875),
    .X(_03840_));
 sky130_fd_sc_hd__nand4_1 _09936_ (.A(net440),
    .B(net932),
    .C(net746),
    .D(net875),
    .Y(_03841_));
 sky130_fd_sc_hd__a22oi_1 _09937_ (.A1(net1393),
    .A2(net1690),
    .B1(_03839_),
    .B2(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__and4_1 _09938_ (.A(net1393),
    .B(net1690),
    .C(_03839_),
    .D(_03841_),
    .X(_03843_));
 sky130_fd_sc_hd__or2_1 _09939_ (.A(_03842_),
    .B(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__nor2_1 _09940_ (.A(_03838_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__o21ai_2 _09941_ (.A1(_03837_),
    .A2(_03845_),
    .B1(_03830_),
    .Y(_03846_));
 sky130_fd_sc_hd__or3_1 _09942_ (.A(_03830_),
    .B(_03837_),
    .C(_03845_),
    .X(_03847_));
 sky130_fd_sc_hd__o211ai_2 _09943_ (.A1(net3683),
    .A2(_03843_),
    .B1(_03846_),
    .C1(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2_1 _09944_ (.A(_03846_),
    .B(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2b_1 _09945_ (.A_N(_03829_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__nor2_1 _09946_ (.A(_03828_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__and2_1 _09947_ (.A(_03828_),
    .B(_03850_),
    .X(_03852_));
 sky130_fd_sc_hd__or2_1 _09948_ (.A(_03851_),
    .B(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__a211o_1 _09949_ (.A1(_03846_),
    .A2(_03847_),
    .B1(net3683),
    .C1(_03843_),
    .X(_03854_));
 sky130_fd_sc_hd__xor2_1 _09950_ (.A(_03838_),
    .B(_03844_),
    .X(_03855_));
 sky130_fd_sc_hd__xnor2_2 _09951_ (.A(_03834_),
    .B(_03835_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand4_2 _09952_ (.A(net812),
    .B(net791),
    .C(net1857),
    .D(net675),
    .Y(_03857_));
 sky130_fd_sc_hd__a22o_1 _09953_ (.A1(net791),
    .A2(net1857),
    .B1(net675),
    .B2(net812),
    .X(_03858_));
 sky130_fd_sc_hd__nand4_2 _09954_ (.A(net863),
    .B(net1870),
    .C(_03857_),
    .D(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(_03857_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__and2b_1 _09956_ (.A_N(_03856_),
    .B(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__xor2_2 _09957_ (.A(_03856_),
    .B(_03860_),
    .X(_03862_));
 sky130_fd_sc_hd__a22o_1 _09958_ (.A1(net2262),
    .A2(net746),
    .B1(net875),
    .B2(net2383),
    .X(_03863_));
 sky130_fd_sc_hd__nand4_1 _09959_ (.A(net3655),
    .B(net2262),
    .C(net746),
    .D(net875),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2_1 _09960_ (.A(_03863_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__nand2_1 _09961_ (.A(net3682),
    .B(net1690),
    .Y(_03866_));
 sky130_fd_sc_hd__xnor2_2 _09962_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__nor2_1 _09963_ (.A(_03862_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__o21a_1 _09964_ (.A1(_03861_),
    .A2(_03868_),
    .B1(_03855_),
    .X(_03869_));
 sky130_fd_sc_hd__or3_1 _09965_ (.A(_03855_),
    .B(_03861_),
    .C(_03868_),
    .X(_03870_));
 sky130_fd_sc_hd__nand2b_1 _09966_ (.A_N(_03869_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__o21ai_2 _09967_ (.A1(_03865_),
    .A2(_03866_),
    .B1(_03864_),
    .Y(_03872_));
 sky130_fd_sc_hd__and2b_1 _09968_ (.A_N(_03871_),
    .B(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__o211ai_4 _09969_ (.A1(_03869_),
    .A2(_03873_),
    .B1(net3684),
    .C1(_03854_),
    .Y(_03874_));
 sky130_fd_sc_hd__xor2_1 _09970_ (.A(_03829_),
    .B(_03849_),
    .X(_03875_));
 sky130_fd_sc_hd__or2_1 _09971_ (.A(_03874_),
    .B(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__a211o_1 _09972_ (.A1(_03848_),
    .A2(_03854_),
    .B1(_03869_),
    .C1(_03873_),
    .X(_03877_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_03874_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_2 _09974_ (.A(_03871_),
    .B(_03872_),
    .Y(_03879_));
 sky130_fd_sc_hd__xor2_2 _09975_ (.A(_03862_),
    .B(_03867_),
    .X(_03880_));
 sky130_fd_sc_hd__a22o_1 _09976_ (.A1(net863),
    .A2(net1870),
    .B1(_03857_),
    .B2(_03858_),
    .X(_03881_));
 sky130_fd_sc_hd__and4_1 _09977_ (.A(net812),
    .B(net791),
    .C(net675),
    .D(net1870),
    .X(_03882_));
 sky130_fd_sc_hd__nand3_1 _09978_ (.A(_03859_),
    .B(_03881_),
    .C(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__a22oi_1 _09979_ (.A1(net1879),
    .A2(net746),
    .B1(net875),
    .B2(net2262),
    .Y(_03884_));
 sky130_fd_sc_hd__and4_1 _09980_ (.A(net2262),
    .B(net1879),
    .C(net2869),
    .D(net875),
    .X(_03885_));
 sky130_fd_sc_hd__nor2_1 _09981_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(net932),
    .B(net1690),
    .Y(_03887_));
 sky130_fd_sc_hd__and3_1 _09983_ (.A(net932),
    .B(net1690),
    .C(_03886_),
    .X(_03888_));
 sky130_fd_sc_hd__xnor2_2 _09984_ (.A(_03886_),
    .B(_03887_),
    .Y(_03889_));
 sky130_fd_sc_hd__a21o_1 _09985_ (.A1(_03859_),
    .A2(_03881_),
    .B1(_03882_),
    .X(_03890_));
 sky130_fd_sc_hd__and3_1 _09986_ (.A(_03883_),
    .B(_03889_),
    .C(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__a21boi_2 _09987_ (.A1(_03889_),
    .A2(_03890_),
    .B1_N(_03883_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2b_1 _09988_ (.A_N(_03892_),
    .B(_03880_),
    .Y(_03893_));
 sky130_fd_sc_hd__xor2_2 _09989_ (.A(_03880_),
    .B(_03892_),
    .X(_03894_));
 sky130_fd_sc_hd__o211a_1 _09990_ (.A1(_03885_),
    .A2(_03888_),
    .B1(net1393),
    .C1(net1767),
    .X(_03895_));
 sky130_fd_sc_hd__a211oi_1 _09991_ (.A1(net1393),
    .A2(net1767),
    .B1(_03885_),
    .C1(_03888_),
    .Y(_03896_));
 sky130_fd_sc_hd__or2_1 _09992_ (.A(_03895_),
    .B(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__o21ai_2 _09993_ (.A1(_03894_),
    .A2(_03897_),
    .B1(_03893_),
    .Y(_03898_));
 sky130_fd_sc_hd__xor2_2 _09994_ (.A(_03879_),
    .B(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__and2_1 _09995_ (.A(_03895_),
    .B(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__a21oi_2 _09996_ (.A1(_03879_),
    .A2(_03898_),
    .B1(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__or2_1 _09997_ (.A(_03878_),
    .B(_03901_),
    .X(_03902_));
 sky130_fd_sc_hd__xnor2_2 _09998_ (.A(_03878_),
    .B(_03901_),
    .Y(_03903_));
 sky130_fd_sc_hd__xnor2_2 _09999_ (.A(_03895_),
    .B(_03899_),
    .Y(_03904_));
 sky130_fd_sc_hd__xnor2_1 _10000_ (.A(_03894_),
    .B(_03897_),
    .Y(_03905_));
 sky130_fd_sc_hd__a21oi_1 _10001_ (.A1(_03883_),
    .A2(_03890_),
    .B1(_03889_),
    .Y(_03906_));
 sky130_fd_sc_hd__a22oi_1 _10002_ (.A1(net791),
    .A2(net675),
    .B1(net1870),
    .B2(net812),
    .Y(_03907_));
 sky130_fd_sc_hd__nor2_1 _10003_ (.A(_03882_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__a22o_1 _10004_ (.A1(net863),
    .A2(net746),
    .B1(net2072),
    .B2(net1879),
    .X(_03909_));
 sky130_fd_sc_hd__nand4_1 _10005_ (.A(net1879),
    .B(net1964),
    .C(net746),
    .D(net2072),
    .Y(_03910_));
 sky130_fd_sc_hd__and2_1 _10006_ (.A(net2262),
    .B(net1690),
    .X(_03911_));
 sky130_fd_sc_hd__a21o_1 _10007_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__nand3_1 _10008_ (.A(_03909_),
    .B(_03910_),
    .C(_03911_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand3_2 _10009_ (.A(_03908_),
    .B(_03912_),
    .C(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__or3_1 _10010_ (.A(_03891_),
    .B(_03906_),
    .C(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a21bo_1 _10011_ (.A1(_03909_),
    .A2(_03911_),
    .B1_N(_03910_),
    .X(_03916_));
 sky130_fd_sc_hd__a21oi_1 _10012_ (.A1(net440),
    .A2(net1767),
    .B1(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__and3_1 _10013_ (.A(net440),
    .B(net1767),
    .C(_03916_),
    .X(_03918_));
 sky130_fd_sc_hd__nor2_1 _10014_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(net1393),
    .B(net821),
    .Y(_03920_));
 sky130_fd_sc_hd__xnor2_1 _10016_ (.A(_03919_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__o21ai_1 _10017_ (.A1(_03891_),
    .A2(_03906_),
    .B1(_03914_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand3_2 _10018_ (.A(_03915_),
    .B(_03921_),
    .C(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_1 _10019_ (.A(_03915_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2b_1 _10020_ (.A_N(_03905_),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__xnor2_1 _10021_ (.A(_03905_),
    .B(_03924_),
    .Y(_03926_));
 sky130_fd_sc_hd__a31o_1 _10022_ (.A1(net1393),
    .A2(net821),
    .A3(_03919_),
    .B1(_03918_),
    .X(_03927_));
 sky130_fd_sc_hd__a21bo_1 _10023_ (.A1(_03926_),
    .A2(_03927_),
    .B1_N(_03925_),
    .X(_03928_));
 sky130_fd_sc_hd__and2b_1 _10024_ (.A_N(_03904_),
    .B(_03928_),
    .X(_03929_));
 sky130_fd_sc_hd__xnor2_2 _10025_ (.A(_03904_),
    .B(_03928_),
    .Y(_03930_));
 sky130_fd_sc_hd__xnor2_1 _10026_ (.A(_03926_),
    .B(_03927_),
    .Y(_03931_));
 sky130_fd_sc_hd__a21o_1 _10027_ (.A1(_03915_),
    .A2(_03922_),
    .B1(_03921_),
    .X(_03932_));
 sky130_fd_sc_hd__a21o_1 _10028_ (.A1(_03912_),
    .A2(_03913_),
    .B1(_03908_),
    .X(_03933_));
 sky130_fd_sc_hd__a22o_1 _10029_ (.A1(net812),
    .A2(net746),
    .B1(net875),
    .B2(net863),
    .X(_03934_));
 sky130_fd_sc_hd__nand4_1 _10030_ (.A(net863),
    .B(net1771),
    .C(net746),
    .D(net875),
    .Y(_03935_));
 sky130_fd_sc_hd__and2_1 _10031_ (.A(net1879),
    .B(net1690),
    .X(_03936_));
 sky130_fd_sc_hd__a21oi_1 _10032_ (.A1(_03934_),
    .A2(_03935_),
    .B1(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__and3_1 _10033_ (.A(_03934_),
    .B(_03935_),
    .C(_03936_),
    .X(_03938_));
 sky130_fd_sc_hd__and4bb_1 _10034_ (.A_N(_03937_),
    .B_N(_03938_),
    .C(net791),
    .D(net1870),
    .X(_03939_));
 sky130_fd_sc_hd__nand3_1 _10035_ (.A(_03914_),
    .B(_03933_),
    .C(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__a21bo_1 _10036_ (.A1(_03934_),
    .A2(_03936_),
    .B1_N(_03935_),
    .X(_03941_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(net932),
    .B(net1767),
    .Y(_03942_));
 sky130_fd_sc_hd__and3_1 _10038_ (.A(net932),
    .B(net1767),
    .C(_03941_),
    .X(_03943_));
 sky130_fd_sc_hd__xnor2_1 _10039_ (.A(_03941_),
    .B(_03942_),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_1 _10040_ (.A(net440),
    .B(net821),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_1 _10041_ (.A(_03944_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__a21o_1 _10042_ (.A1(_03914_),
    .A2(_03933_),
    .B1(_03939_),
    .X(_03947_));
 sky130_fd_sc_hd__nand3_1 _10043_ (.A(_03940_),
    .B(_03946_),
    .C(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(_03940_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__nand3_1 _10045_ (.A(_03923_),
    .B(_03932_),
    .C(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__a31o_1 _10046_ (.A1(net440),
    .A2(net821),
    .A3(_03944_),
    .B1(_03943_),
    .X(_03951_));
 sky130_fd_sc_hd__a21o_1 _10047_ (.A1(_03923_),
    .A2(_03932_),
    .B1(_03949_),
    .X(_03952_));
 sky130_fd_sc_hd__and3_1 _10048_ (.A(_03950_),
    .B(_03951_),
    .C(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__a31o_1 _10049_ (.A1(_03923_),
    .A2(_03932_),
    .A3(_03949_),
    .B1(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__and2b_1 _10050_ (.A_N(_03931_),
    .B(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__xnor2_1 _10051_ (.A(_03931_),
    .B(_03954_),
    .Y(_03956_));
 sky130_fd_sc_hd__a21oi_1 _10052_ (.A1(_03950_),
    .A2(_03952_),
    .B1(_03951_),
    .Y(_03957_));
 sky130_fd_sc_hd__a21o_1 _10053_ (.A1(_03940_),
    .A2(_03947_),
    .B1(_03946_),
    .X(_03958_));
 sky130_fd_sc_hd__o2bb2a_1 _10054_ (.A1_N(net791),
    .A2_N(net1870),
    .B1(_03937_),
    .B2(_03938_),
    .X(_03959_));
 sky130_fd_sc_hd__nor2_1 _10055_ (.A(_03939_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _10056_ (.A(net932),
    .B(net821),
    .Y(_03961_));
 sky130_fd_sc_hd__and3_1 _10057_ (.A(net812),
    .B(net791),
    .C(net875),
    .X(_03962_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(net863),
    .B(net1690),
    .Y(_03963_));
 sky130_fd_sc_hd__a22o_1 _10059_ (.A1(net791),
    .A2(net746),
    .B1(net875),
    .B2(net812),
    .X(_03964_));
 sky130_fd_sc_hd__a21bo_1 _10060_ (.A1(net746),
    .A2(_03962_),
    .B1_N(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__a32o_1 _10061_ (.A1(net863),
    .A2(net1690),
    .A3(_03964_),
    .B1(_03962_),
    .B2(net746),
    .X(_03966_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(net2262),
    .B(net1767),
    .Y(_03967_));
 sky130_fd_sc_hd__and3_1 _10063_ (.A(net2262),
    .B(net1767),
    .C(_03966_),
    .X(_03968_));
 sky130_fd_sc_hd__xnor2_1 _10064_ (.A(_03966_),
    .B(_03967_),
    .Y(_03969_));
 sky130_fd_sc_hd__xnor2_1 _10065_ (.A(_03961_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__and2_1 _10066_ (.A(_03960_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nand3_2 _10067_ (.A(_03948_),
    .B(_03958_),
    .C(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__a31o_1 _10068_ (.A1(net932),
    .A2(net821),
    .A3(_03969_),
    .B1(_03968_),
    .X(_03973_));
 sky130_fd_sc_hd__a21o_1 _10069_ (.A1(_03948_),
    .A2(_03958_),
    .B1(_03971_),
    .X(_03974_));
 sky130_fd_sc_hd__nand3_2 _10070_ (.A(_03972_),
    .B(_03973_),
    .C(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__a211oi_1 _10071_ (.A1(_03972_),
    .A2(_03975_),
    .B1(_03953_),
    .C1(_03957_),
    .Y(_03976_));
 sky130_fd_sc_hd__o211ai_2 _10072_ (.A1(_03953_),
    .A2(_03957_),
    .B1(_03972_),
    .C1(_03975_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2b_1 _10073_ (.A_N(_03976_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a21o_1 _10074_ (.A1(_03972_),
    .A2(_03974_),
    .B1(_03973_),
    .X(_03979_));
 sky130_fd_sc_hd__xnor2_1 _10075_ (.A(_03960_),
    .B(_03970_),
    .Y(_03980_));
 sky130_fd_sc_hd__xor2_1 _10076_ (.A(_03963_),
    .B(_03965_),
    .X(_03981_));
 sky130_fd_sc_hd__and4_1 _10077_ (.A(net812),
    .B(net791),
    .C(net875),
    .D(net1690),
    .X(_03982_));
 sky130_fd_sc_hd__inv_2 _10078_ (.A(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(net1879),
    .B(net1767),
    .Y(_03984_));
 sky130_fd_sc_hd__nor2_1 _10080_ (.A(_03983_),
    .B(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__xnor2_1 _10081_ (.A(_03982_),
    .B(_03984_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _10082_ (.A(net2262),
    .B(net821),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_1 _10083_ (.A(_03986_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_1 _10084_ (.A(_03981_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__nor2_1 _10085_ (.A(_03980_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__a31o_1 _10086_ (.A1(net2262),
    .A2(net821),
    .A3(_03986_),
    .B1(_03985_),
    .X(_03991_));
 sky130_fd_sc_hd__xor2_1 _10087_ (.A(_03980_),
    .B(_03989_),
    .X(_03992_));
 sky130_fd_sc_hd__a21o_1 _10088_ (.A1(_03991_),
    .A2(_03992_),
    .B1(_03990_),
    .X(_03993_));
 sky130_fd_sc_hd__and3_1 _10089_ (.A(_03975_),
    .B(_03979_),
    .C(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__a21o_1 _10090_ (.A1(_03975_),
    .A2(_03979_),
    .B1(_03993_),
    .X(_03995_));
 sky130_fd_sc_hd__and2b_1 _10091_ (.A_N(_03994_),
    .B(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__xnor2_1 _10092_ (.A(_03991_),
    .B(_03992_),
    .Y(_03997_));
 sky130_fd_sc_hd__xnor2_1 _10093_ (.A(_03981_),
    .B(_03988_),
    .Y(_03998_));
 sky130_fd_sc_hd__and4_1 _10094_ (.A(net1879),
    .B(net863),
    .C(net1767),
    .D(net821),
    .X(_03999_));
 sky130_fd_sc_hd__inv_2 _10095_ (.A(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__a22o_1 _10096_ (.A1(net791),
    .A2(net875),
    .B1(net1690),
    .B2(net812),
    .X(_04001_));
 sky130_fd_sc_hd__a22o_1 _10097_ (.A1(net863),
    .A2(net1767),
    .B1(net821),
    .B2(net1879),
    .X(_04002_));
 sky130_fd_sc_hd__or4bb_2 _10098_ (.A(_03982_),
    .B(_03999_),
    .C_N(_04001_),
    .D_N(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__a21o_1 _10099_ (.A1(_04000_),
    .A2(_04003_),
    .B1(_03998_),
    .X(_04004_));
 sky130_fd_sc_hd__nand3_1 _10100_ (.A(_03998_),
    .B(_04000_),
    .C(_04003_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_04004_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__a22o_1 _10102_ (.A1(_03983_),
    .A2(_04001_),
    .B1(_04002_),
    .B2(_04000_),
    .X(_04007_));
 sky130_fd_sc_hd__and4_1 _10103_ (.A(net863),
    .B(net812),
    .C(net1767),
    .D(net821),
    .X(_04008_));
 sky130_fd_sc_hd__a22o_1 _10104_ (.A1(net812),
    .A2(net1767),
    .B1(net2808),
    .B2(net863),
    .X(_04009_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__and4b_1 _10106_ (.A_N(_04008_),
    .B(_04009_),
    .C(net791),
    .D(net1690),
    .X(_04011_));
 sky130_fd_sc_hd__or2_1 _10107_ (.A(_04008_),
    .B(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__and3_1 _10108_ (.A(_04003_),
    .B(_04007_),
    .C(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__o2bb2a_1 _10109_ (.A1_N(net1630),
    .A2_N(net1690),
    .B1(_04008_),
    .B2(_04010_),
    .X(_04014_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04011_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__and4_1 _10111_ (.A(net1773),
    .B(net1632),
    .C(net1767),
    .D(net821),
    .X(_04016_));
 sky130_fd_sc_hd__and2_2 _10112_ (.A(_04015_),
    .B(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__a21oi_1 _10113_ (.A1(_04003_),
    .A2(_04007_),
    .B1(_04012_),
    .Y(_04018_));
 sky130_fd_sc_hd__nor2_1 _10114_ (.A(_04013_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__a21oi_2 _10115_ (.A1(_04017_),
    .A2(_04019_),
    .B1(_04013_),
    .Y(_04020_));
 sky130_fd_sc_hd__or2_1 _10116_ (.A(_04006_),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__a21oi_2 _10117_ (.A1(_04004_),
    .A2(_04021_),
    .B1(_03997_),
    .Y(_04022_));
 sky130_fd_sc_hd__a21o_1 _10118_ (.A1(_03995_),
    .A2(_04022_),
    .B1(_03994_),
    .X(_04023_));
 sky130_fd_sc_hd__a21o_1 _10119_ (.A1(_03977_),
    .A2(_04023_),
    .B1(_03976_),
    .X(_04024_));
 sky130_fd_sc_hd__and2_1 _10120_ (.A(_03956_),
    .B(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__a21o_1 _10121_ (.A1(_03956_),
    .A2(_04024_),
    .B1(_03955_),
    .X(_04026_));
 sky130_fd_sc_hd__a21oi_2 _10122_ (.A1(_03930_),
    .A2(_04026_),
    .B1(_03929_),
    .Y(_04027_));
 sky130_fd_sc_hd__o21ai_1 _10123_ (.A1(_03903_),
    .A2(_04027_),
    .B1(_03902_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2b_1 _10124_ (.A_N(_03875_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__a21oi_1 _10125_ (.A1(_03876_),
    .A2(_04029_),
    .B1(_03853_),
    .Y(_04030_));
 sky130_fd_sc_hd__and3_1 _10126_ (.A(_03853_),
    .B(_03876_),
    .C(_04029_),
    .X(_04031_));
 sky130_fd_sc_hd__or2_1 _10127_ (.A(_04030_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__xnor2_1 _10128_ (.A(_03527_),
    .B(_03780_),
    .Y(_04033_));
 sky130_fd_sc_hd__or2_1 _10129_ (.A(_04032_),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(net2792),
    .B(net2315),
    .Y(_04035_));
 sky130_fd_sc_hd__a22o_1 _10131_ (.A1(net854),
    .A2(net1930),
    .B1(net707),
    .B2(net473),
    .X(_04036_));
 sky130_fd_sc_hd__and3_1 _10132_ (.A(net473),
    .B(net1930),
    .C(net707),
    .X(_04037_));
 sky130_fd_sc_hd__a21bo_1 _10133_ (.A1(net854),
    .A2(_04037_),
    .B1_N(_04036_),
    .X(_04038_));
 sky130_fd_sc_hd__nand2_1 _10134_ (.A(net1429),
    .B(net1938),
    .Y(_04039_));
 sky130_fd_sc_hd__xnor2_1 _10135_ (.A(_04038_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__and4_1 _10136_ (.A(net854),
    .B(net2101),
    .C(net1930),
    .D(net707),
    .X(_04041_));
 sky130_fd_sc_hd__a22o_1 _10137_ (.A1(net2101),
    .A2(net1930),
    .B1(net707),
    .B2(net854),
    .X(_04042_));
 sky130_fd_sc_hd__inv_2 _10138_ (.A(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__and4b_1 _10139_ (.A_N(_04041_),
    .B(_04042_),
    .C(net473),
    .D(net1938),
    .X(_04044_));
 sky130_fd_sc_hd__nor2_1 _10140_ (.A(_04041_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__or2_1 _10141_ (.A(_04040_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__xnor2_1 _10142_ (.A(_04040_),
    .B(_04045_),
    .Y(_04047_));
 sky130_fd_sc_hd__o2bb2a_1 _10143_ (.A1_N(net473),
    .A2_N(net1938),
    .B1(_04041_),
    .B2(_04043_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _10144_ (.A(_04044_),
    .B(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__nand4_1 _10145_ (.A(net2101),
    .B(net1825),
    .C(net1930),
    .D(net707),
    .Y(_04050_));
 sky130_fd_sc_hd__a22o_1 _10146_ (.A1(net1825),
    .A2(net1930),
    .B1(net707),
    .B2(net2101),
    .X(_04051_));
 sky130_fd_sc_hd__nand2_1 _10147_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_1 _10148_ (.A(net854),
    .B(net1938),
    .Y(_04053_));
 sky130_fd_sc_hd__o21ai_1 _10149_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04050_),
    .Y(_04054_));
 sky130_fd_sc_hd__and2b_1 _10150_ (.A_N(_04049_),
    .B(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__and2b_1 _10151_ (.A_N(_04054_),
    .B(_04049_),
    .X(_04056_));
 sky130_fd_sc_hd__nor2_1 _10152_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(net1429),
    .B(net794),
    .Y(_04058_));
 sky130_fd_sc_hd__a31oi_1 _10154_ (.A1(net1429),
    .A2(net794),
    .A3(_04057_),
    .B1(_04055_),
    .Y(_04059_));
 sky130_fd_sc_hd__or2_1 _10155_ (.A(_04047_),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__nand2_1 _10156_ (.A(_04047_),
    .B(_04059_),
    .Y(_04061_));
 sky130_fd_sc_hd__and2_1 _10157_ (.A(_04060_),
    .B(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__xnor2_1 _10158_ (.A(_04057_),
    .B(_04058_),
    .Y(_04063_));
 sky130_fd_sc_hd__xnor2_1 _10159_ (.A(_04052_),
    .B(_04053_),
    .Y(_04064_));
 sky130_fd_sc_hd__and4_1 _10160_ (.A(net1825),
    .B(net43),
    .C(net1930),
    .D(net707),
    .X(_04065_));
 sky130_fd_sc_hd__a22oi_1 _10161_ (.A1(net43),
    .A2(net1930),
    .B1(net707),
    .B2(net1825),
    .Y(_04066_));
 sky130_fd_sc_hd__or2_1 _10162_ (.A(_04065_),
    .B(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__nand2_1 _10163_ (.A(net2101),
    .B(net1938),
    .Y(_04068_));
 sky130_fd_sc_hd__o21ba_1 _10164_ (.A1(_04067_),
    .A2(_04068_),
    .B1_N(_04065_),
    .X(_04069_));
 sky130_fd_sc_hd__xnor2_1 _10165_ (.A(_04064_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__a22oi_2 _10166_ (.A1(net473),
    .A2(net794),
    .B1(net869),
    .B2(net1429),
    .Y(_04071_));
 sky130_fd_sc_hd__and4_1 _10167_ (.A(net1429),
    .B(net473),
    .C(net2475),
    .D(net869),
    .X(_04072_));
 sky130_fd_sc_hd__nor2_1 _10168_ (.A(_04071_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__o32a_1 _10169_ (.A1(_04070_),
    .A2(_04071_),
    .A3(_04072_),
    .B1(_04069_),
    .B2(_04064_),
    .X(_04074_));
 sky130_fd_sc_hd__and2b_1 _10170_ (.A_N(_04074_),
    .B(_04063_),
    .X(_04075_));
 sky130_fd_sc_hd__xnor2_1 _10171_ (.A(_04063_),
    .B(_04074_),
    .Y(_04076_));
 sky130_fd_sc_hd__a21oi_1 _10172_ (.A1(_04072_),
    .A2(_04076_),
    .B1(_04075_),
    .Y(_04077_));
 sky130_fd_sc_hd__and2b_1 _10173_ (.A_N(_04077_),
    .B(_04062_),
    .X(_04078_));
 sky130_fd_sc_hd__a22oi_1 _10174_ (.A1(net2792),
    .A2(net1930),
    .B1(net707),
    .B2(net1429),
    .Y(_04079_));
 sky130_fd_sc_hd__and4_1 _10175_ (.A(net1429),
    .B(net2792),
    .C(net1930),
    .D(net2315),
    .X(_04080_));
 sky130_fd_sc_hd__nor2_1 _10176_ (.A(_04079_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a32o_1 _10177_ (.A1(net1429),
    .A2(net1938),
    .A3(_04036_),
    .B1(_04037_),
    .B2(net854),
    .X(_04082_));
 sky130_fd_sc_hd__nand2_1 _10178_ (.A(_04081_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__or2_1 _10179_ (.A(_04081_),
    .B(_04082_),
    .X(_04084_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _10181_ (.A(_04046_),
    .B(_04060_),
    .Y(_04086_));
 sky130_fd_sc_hd__xnor2_1 _10182_ (.A(_04085_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(_04078_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__or2_1 _10184_ (.A(_04078_),
    .B(_04087_),
    .X(_04089_));
 sky130_fd_sc_hd__and2_1 _10185_ (.A(_04088_),
    .B(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__inv_2 _10186_ (.A(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__and2b_1 _10187_ (.A_N(_04062_),
    .B(_04077_),
    .X(_04092_));
 sky130_fd_sc_hd__or2_1 _10188_ (.A(_04078_),
    .B(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__xnor2_1 _10189_ (.A(_04072_),
    .B(_04076_),
    .Y(_04094_));
 sky130_fd_sc_hd__xnor2_1 _10190_ (.A(_04070_),
    .B(_04073_),
    .Y(_04095_));
 sky130_fd_sc_hd__xnor2_1 _10191_ (.A(_04067_),
    .B(_04068_),
    .Y(_04096_));
 sky130_fd_sc_hd__and4_1 _10192_ (.A(net43),
    .B(net914),
    .C(net1930),
    .D(net707),
    .X(_04097_));
 sky130_fd_sc_hd__a22o_1 _10193_ (.A1(net914),
    .A2(net1930),
    .B1(net707),
    .B2(net43),
    .X(_04098_));
 sky130_fd_sc_hd__nand2b_1 _10194_ (.A_N(_04097_),
    .B(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(net1825),
    .B(net1938),
    .Y(_04100_));
 sky130_fd_sc_hd__a31o_1 _10196_ (.A1(net1825),
    .A2(net1938),
    .A3(_04098_),
    .B1(_04097_),
    .X(_04101_));
 sky130_fd_sc_hd__and2b_1 _10197_ (.A_N(_04096_),
    .B(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__xor2_1 _10198_ (.A(_04096_),
    .B(_04101_),
    .X(_04103_));
 sky130_fd_sc_hd__a22o_1 _10199_ (.A1(net854),
    .A2(net794),
    .B1(net869),
    .B2(net473),
    .X(_04104_));
 sky130_fd_sc_hd__and4_1 _10200_ (.A(net473),
    .B(net854),
    .C(net2475),
    .D(net869),
    .X(_04105_));
 sky130_fd_sc_hd__nand4_1 _10201_ (.A(net473),
    .B(net2453),
    .C(net794),
    .D(net869),
    .Y(_04106_));
 sky130_fd_sc_hd__a22oi_1 _10202_ (.A1(net1429),
    .A2(net1717),
    .B1(_04104_),
    .B2(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__and4_1 _10203_ (.A(net1429),
    .B(net1717),
    .C(_04104_),
    .D(_04106_),
    .X(_04108_));
 sky130_fd_sc_hd__or2_1 _10204_ (.A(_04107_),
    .B(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(_04103_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__o21ai_1 _10206_ (.A1(_04102_),
    .A2(_04110_),
    .B1(_04095_),
    .Y(_04111_));
 sky130_fd_sc_hd__or3_1 _10207_ (.A(_04095_),
    .B(_04102_),
    .C(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _10208_ (.A(_04111_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nor2_1 _10209_ (.A(_04105_),
    .B(_04108_),
    .Y(_04114_));
 sky130_fd_sc_hd__or2_1 _10210_ (.A(_04113_),
    .B(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a21o_1 _10211_ (.A1(_04111_),
    .A2(_04115_),
    .B1(_04094_),
    .X(_04116_));
 sky130_fd_sc_hd__or2_1 _10212_ (.A(_04093_),
    .B(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(_04093_),
    .B(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__and2_1 _10214_ (.A(_04117_),
    .B(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__inv_2 _10215_ (.A(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__nand3_1 _10216_ (.A(_04094_),
    .B(_04111_),
    .C(_04115_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _10217_ (.A(_04116_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__xnor2_1 _10218_ (.A(_04113_),
    .B(_04114_),
    .Y(_04123_));
 sky130_fd_sc_hd__xor2_1 _10219_ (.A(_04103_),
    .B(_04109_),
    .X(_04124_));
 sky130_fd_sc_hd__xnor2_1 _10220_ (.A(_04099_),
    .B(_04100_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand4_2 _10221_ (.A(net914),
    .B(net731),
    .C(net1930),
    .D(net707),
    .Y(_04126_));
 sky130_fd_sc_hd__a22o_1 _10222_ (.A1(net731),
    .A2(net1930),
    .B1(net707),
    .B2(net914),
    .X(_04127_));
 sky130_fd_sc_hd__nand4_2 _10223_ (.A(net43),
    .B(net1938),
    .C(_04126_),
    .D(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__nand2_1 _10224_ (.A(_04126_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__and2b_1 _10225_ (.A_N(_04125_),
    .B(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__xor2_1 _10226_ (.A(_04125_),
    .B(_04129_),
    .X(_04131_));
 sky130_fd_sc_hd__a22o_1 _10227_ (.A1(net2101),
    .A2(net794),
    .B1(net869),
    .B2(net854),
    .X(_04132_));
 sky130_fd_sc_hd__nand4_2 _10228_ (.A(net854),
    .B(net2101),
    .C(net2475),
    .D(net869),
    .Y(_04133_));
 sky130_fd_sc_hd__a22o_1 _10229_ (.A1(net473),
    .A2(net1717),
    .B1(_04132_),
    .B2(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__nand4_2 _10230_ (.A(net473),
    .B(net1717),
    .C(_04132_),
    .D(_04133_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand2_1 _10231_ (.A(_04134_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_1 _10232_ (.A(_04131_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__o21a_1 _10233_ (.A1(_04130_),
    .A2(_04137_),
    .B1(_04124_),
    .X(_04138_));
 sky130_fd_sc_hd__nor3_1 _10234_ (.A(_04124_),
    .B(_04130_),
    .C(_04137_),
    .Y(_04139_));
 sky130_fd_sc_hd__a211oi_1 _10235_ (.A1(_04133_),
    .A2(_04135_),
    .B1(_04138_),
    .C1(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__or2_1 _10236_ (.A(_04138_),
    .B(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__nand2b_1 _10237_ (.A_N(_04123_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__xor2_1 _10238_ (.A(_04122_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__xnor2_1 _10239_ (.A(_04123_),
    .B(_04141_),
    .Y(_04144_));
 sky130_fd_sc_hd__o211ai_1 _10240_ (.A1(_04138_),
    .A2(_04139_),
    .B1(_04133_),
    .C1(_04135_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2b_1 _10241_ (.A_N(_04140_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__xor2_1 _10242_ (.A(_04131_),
    .B(_04136_),
    .X(_04147_));
 sky130_fd_sc_hd__a22o_1 _10243_ (.A1(net43),
    .A2(net1938),
    .B1(_04126_),
    .B2(_04127_),
    .X(_04148_));
 sky130_fd_sc_hd__and4_1 _10244_ (.A(net914),
    .B(net731),
    .C(net707),
    .D(net1938),
    .X(_04149_));
 sky130_fd_sc_hd__and3_1 _10245_ (.A(_04128_),
    .B(_04148_),
    .C(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__nand3_1 _10246_ (.A(_04128_),
    .B(_04148_),
    .C(_04149_),
    .Y(_04151_));
 sky130_fd_sc_hd__a21o_1 _10247_ (.A1(_04128_),
    .A2(_04148_),
    .B1(_04149_),
    .X(_04152_));
 sky130_fd_sc_hd__a22oi_2 _10248_ (.A1(net1825),
    .A2(net794),
    .B1(net2481),
    .B2(net2101),
    .Y(_04153_));
 sky130_fd_sc_hd__and4_1 _10249_ (.A(net2101),
    .B(net1825),
    .C(net794),
    .D(net2481),
    .X(_04154_));
 sky130_fd_sc_hd__nor2_1 _10250_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(net854),
    .B(net1717),
    .Y(_04156_));
 sky130_fd_sc_hd__xnor2_1 _10252_ (.A(_04155_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__and3_1 _10253_ (.A(_04151_),
    .B(_04152_),
    .C(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__o21a_1 _10254_ (.A1(_04150_),
    .A2(_04158_),
    .B1(_04147_),
    .X(_04159_));
 sky130_fd_sc_hd__nor3_1 _10255_ (.A(_04147_),
    .B(_04150_),
    .C(_04158_),
    .Y(_04160_));
 sky130_fd_sc_hd__o21ba_1 _10256_ (.A1(_04153_),
    .A2(_04156_),
    .B1_N(_04154_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _10257_ (.A(net1429),
    .B(net1713),
    .Y(_04162_));
 sky130_fd_sc_hd__nor2_1 _10258_ (.A(_04161_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__xnor2_1 _10259_ (.A(_04161_),
    .B(_04162_),
    .Y(_04164_));
 sky130_fd_sc_hd__nor3_1 _10260_ (.A(_04159_),
    .B(_04160_),
    .C(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__or2_1 _10261_ (.A(_04159_),
    .B(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__and2b_1 _10262_ (.A_N(_04146_),
    .B(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__xnor2_1 _10263_ (.A(_04146_),
    .B(_04166_),
    .Y(_04168_));
 sky130_fd_sc_hd__and2_1 _10264_ (.A(_04163_),
    .B(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__o21a_1 _10265_ (.A1(_04167_),
    .A2(_04169_),
    .B1(_04144_),
    .X(_04170_));
 sky130_fd_sc_hd__nor3_1 _10266_ (.A(_04144_),
    .B(_04167_),
    .C(_04169_),
    .Y(_04171_));
 sky130_fd_sc_hd__or2_1 _10267_ (.A(_04170_),
    .B(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__xnor2_1 _10268_ (.A(_04163_),
    .B(_04168_),
    .Y(_04173_));
 sky130_fd_sc_hd__o21a_1 _10269_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_04164_),
    .X(_04174_));
 sky130_fd_sc_hd__a21oi_1 _10270_ (.A1(_04151_),
    .A2(_04152_),
    .B1(_04157_),
    .Y(_04175_));
 sky130_fd_sc_hd__a22oi_1 _10271_ (.A1(net731),
    .A2(net707),
    .B1(net1938),
    .B2(net3447),
    .Y(_04176_));
 sky130_fd_sc_hd__nor2_1 _10272_ (.A(_04149_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__a22o_1 _10273_ (.A1(net43),
    .A2(net794),
    .B1(net869),
    .B2(net1825),
    .X(_04178_));
 sky130_fd_sc_hd__nand4_2 _10274_ (.A(net1825),
    .B(net43),
    .C(net794),
    .D(net869),
    .Y(_04179_));
 sky130_fd_sc_hd__and2_1 _10275_ (.A(net2101),
    .B(net1717),
    .X(_04180_));
 sky130_fd_sc_hd__a21o_1 _10276_ (.A1(_04178_),
    .A2(_04179_),
    .B1(_04180_),
    .X(_04181_));
 sky130_fd_sc_hd__nand3_1 _10277_ (.A(_04178_),
    .B(_04179_),
    .C(_04180_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand3_1 _10278_ (.A(_04177_),
    .B(_04181_),
    .C(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__or3_2 _10279_ (.A(_04158_),
    .B(_04175_),
    .C(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__o21ai_1 _10280_ (.A1(_04158_),
    .A2(_04175_),
    .B1(_04183_),
    .Y(_04185_));
 sky130_fd_sc_hd__a21bo_1 _10281_ (.A1(_04178_),
    .A2(_04180_),
    .B1_N(_04179_),
    .X(_04186_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(net473),
    .B(net1713),
    .Y(_04187_));
 sky130_fd_sc_hd__and3_1 _10283_ (.A(net473),
    .B(net1713),
    .C(_04186_),
    .X(_04188_));
 sky130_fd_sc_hd__xnor2_1 _10284_ (.A(_04186_),
    .B(_04187_),
    .Y(_04189_));
 sky130_fd_sc_hd__and2_1 _10285_ (.A(net1429),
    .B(net1926),
    .X(_04190_));
 sky130_fd_sc_hd__nor2_1 _10286_ (.A(_04189_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__and2_1 _10287_ (.A(_04189_),
    .B(_04190_),
    .X(_04192_));
 sky130_fd_sc_hd__nor2_1 _10288_ (.A(_04191_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__nand3_2 _10289_ (.A(_04184_),
    .B(_04185_),
    .C(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__a211o_1 _10290_ (.A1(_04184_),
    .A2(_04194_),
    .B1(_04165_),
    .C1(_04174_),
    .X(_04195_));
 sky130_fd_sc_hd__o211ai_2 _10291_ (.A1(_04165_),
    .A2(_04174_),
    .B1(_04184_),
    .C1(_04194_),
    .Y(_04196_));
 sky130_fd_sc_hd__o211ai_2 _10292_ (.A1(_04188_),
    .A2(_04192_),
    .B1(_04195_),
    .C1(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__nand2b_1 _10294_ (.A_N(_04173_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__xnor2_1 _10295_ (.A(_04173_),
    .B(_04198_),
    .Y(_04200_));
 sky130_fd_sc_hd__a211o_1 _10296_ (.A1(_04195_),
    .A2(_04196_),
    .B1(_04188_),
    .C1(_04192_),
    .X(_04201_));
 sky130_fd_sc_hd__a21o_1 _10297_ (.A1(_04184_),
    .A2(_04185_),
    .B1(_04193_),
    .X(_04202_));
 sky130_fd_sc_hd__a21o_1 _10298_ (.A1(_04181_),
    .A2(_04182_),
    .B1(_04177_),
    .X(_04203_));
 sky130_fd_sc_hd__a22o_1 _10299_ (.A1(net914),
    .A2(net794),
    .B1(net869),
    .B2(net43),
    .X(_04204_));
 sky130_fd_sc_hd__nand4_1 _10300_ (.A(net43),
    .B(net914),
    .C(net794),
    .D(net869),
    .Y(_04205_));
 sky130_fd_sc_hd__and2_1 _10301_ (.A(net1825),
    .B(net1717),
    .X(_04206_));
 sky130_fd_sc_hd__a21oi_1 _10302_ (.A1(_04204_),
    .A2(_04205_),
    .B1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__and3_1 _10303_ (.A(_04204_),
    .B(_04205_),
    .C(_04206_),
    .X(_04208_));
 sky130_fd_sc_hd__and4bb_1 _10304_ (.A_N(_04207_),
    .B_N(_04208_),
    .C(net731),
    .D(net1938),
    .X(_04209_));
 sky130_fd_sc_hd__nand3_1 _10305_ (.A(_04183_),
    .B(_04203_),
    .C(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__a21o_1 _10306_ (.A1(_04183_),
    .A2(_04203_),
    .B1(_04209_),
    .X(_04211_));
 sky130_fd_sc_hd__a21bo_1 _10307_ (.A1(_04204_),
    .A2(_04206_),
    .B1_N(_04205_),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_1 _10308_ (.A(net2455),
    .B(net1713),
    .Y(_04213_));
 sky130_fd_sc_hd__and3_1 _10309_ (.A(net2455),
    .B(net1713),
    .C(_04212_),
    .X(_04214_));
 sky130_fd_sc_hd__xnor2_1 _10310_ (.A(_04212_),
    .B(_04213_),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(net473),
    .B(net1926),
    .Y(_04216_));
 sky130_fd_sc_hd__and3_1 _10312_ (.A(net473),
    .B(net1926),
    .C(_04215_),
    .X(_04217_));
 sky130_fd_sc_hd__xnor2_1 _10313_ (.A(_04215_),
    .B(_04216_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand3_1 _10314_ (.A(_04210_),
    .B(_04211_),
    .C(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_1 _10315_ (.A(_04210_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand3_1 _10316_ (.A(_04194_),
    .B(_04202_),
    .C(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a21o_1 _10317_ (.A1(_04194_),
    .A2(_04202_),
    .B1(_04220_),
    .X(_04222_));
 sky130_fd_sc_hd__o211a_1 _10318_ (.A1(_04214_),
    .A2(_04217_),
    .B1(_04221_),
    .C1(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__a31o_1 _10319_ (.A1(_04194_),
    .A2(_04202_),
    .A3(_04220_),
    .B1(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__and3_1 _10320_ (.A(_04197_),
    .B(_04201_),
    .C(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__a21oi_1 _10321_ (.A1(_04197_),
    .A2(_04201_),
    .B1(_04224_),
    .Y(_04226_));
 sky130_fd_sc_hd__a211oi_2 _10322_ (.A1(_04221_),
    .A2(_04222_),
    .B1(_04214_),
    .C1(_04217_),
    .Y(_04227_));
 sky130_fd_sc_hd__o2bb2a_1 _10323_ (.A1_N(net3205),
    .A2_N(net1938),
    .B1(_04207_),
    .B2(_04208_),
    .X(_04228_));
 sky130_fd_sc_hd__nor2_1 _10324_ (.A(_04209_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__and3_1 _10325_ (.A(net914),
    .B(net731),
    .C(net869),
    .X(_04230_));
 sky130_fd_sc_hd__nand2_1 _10326_ (.A(net43),
    .B(net1717),
    .Y(_04231_));
 sky130_fd_sc_hd__a22o_1 _10327_ (.A1(net731),
    .A2(net794),
    .B1(net869),
    .B2(net914),
    .X(_04232_));
 sky130_fd_sc_hd__a21bo_1 _10328_ (.A1(net794),
    .A2(_04230_),
    .B1_N(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__a32o_1 _10329_ (.A1(net43),
    .A2(net1717),
    .A3(_04232_),
    .B1(_04230_),
    .B2(net794),
    .X(_04234_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(net2101),
    .B(net1713),
    .Y(_04235_));
 sky130_fd_sc_hd__and3_1 _10331_ (.A(net2101),
    .B(net1713),
    .C(_04234_),
    .X(_04236_));
 sky130_fd_sc_hd__xnor2_1 _10332_ (.A(_04234_),
    .B(_04235_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(net2455),
    .B(net1926),
    .Y(_04238_));
 sky130_fd_sc_hd__xnor2_1 _10334_ (.A(_04237_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__and2_1 _10335_ (.A(_04229_),
    .B(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__a21o_1 _10336_ (.A1(_04210_),
    .A2(_04211_),
    .B1(_04218_),
    .X(_04241_));
 sky130_fd_sc_hd__nand3_2 _10337_ (.A(_04219_),
    .B(_04240_),
    .C(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__a31o_1 _10338_ (.A1(net2455),
    .A2(net1926),
    .A3(_04237_),
    .B1(_04236_),
    .X(_04243_));
 sky130_fd_sc_hd__a21o_1 _10339_ (.A1(_04219_),
    .A2(_04241_),
    .B1(_04240_),
    .X(_04244_));
 sky130_fd_sc_hd__nand3_2 _10340_ (.A(_04242_),
    .B(_04243_),
    .C(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__a211oi_2 _10341_ (.A1(_04242_),
    .A2(_04245_),
    .B1(_04223_),
    .C1(_04227_),
    .Y(_04246_));
 sky130_fd_sc_hd__inv_2 _10342_ (.A(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__o211a_1 _10343_ (.A1(_04223_),
    .A2(_04227_),
    .B1(_04242_),
    .C1(_04245_),
    .X(_04248_));
 sky130_fd_sc_hd__a21o_1 _10344_ (.A1(_04242_),
    .A2(_04244_),
    .B1(_04243_),
    .X(_04249_));
 sky130_fd_sc_hd__xor2_1 _10345_ (.A(_04231_),
    .B(_04233_),
    .X(_04250_));
 sky130_fd_sc_hd__and4_1 _10346_ (.A(net914),
    .B(net731),
    .C(net869),
    .D(net1717),
    .X(_04251_));
 sky130_fd_sc_hd__inv_2 _10347_ (.A(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _10348_ (.A(net1825),
    .B(net1713),
    .Y(_04253_));
 sky130_fd_sc_hd__nor2_1 _10349_ (.A(_04252_),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__xnor2_1 _10350_ (.A(_04251_),
    .B(_04253_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_1 _10351_ (.A(net2101),
    .B(net1926),
    .Y(_04256_));
 sky130_fd_sc_hd__xnor2_1 _10352_ (.A(_04255_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _10353_ (.A(_04250_),
    .B(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__xnor2_1 _10354_ (.A(_04229_),
    .B(_04239_),
    .Y(_04259_));
 sky130_fd_sc_hd__nor2_1 _10355_ (.A(_04258_),
    .B(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__a31o_1 _10356_ (.A1(net2101),
    .A2(net1926),
    .A3(_04255_),
    .B1(_04254_),
    .X(_04261_));
 sky130_fd_sc_hd__xor2_1 _10357_ (.A(_04258_),
    .B(_04259_),
    .X(_04262_));
 sky130_fd_sc_hd__a21o_1 _10358_ (.A1(_04261_),
    .A2(_04262_),
    .B1(_04260_),
    .X(_04263_));
 sky130_fd_sc_hd__and3_1 _10359_ (.A(_04245_),
    .B(_04249_),
    .C(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__nand3_1 _10360_ (.A(_04245_),
    .B(_04249_),
    .C(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__a21oi_1 _10361_ (.A1(_04245_),
    .A2(_04249_),
    .B1(_04263_),
    .Y(_04266_));
 sky130_fd_sc_hd__xnor2_1 _10362_ (.A(_04261_),
    .B(_04262_),
    .Y(_04267_));
 sky130_fd_sc_hd__xnor2_1 _10363_ (.A(_04250_),
    .B(_04257_),
    .Y(_04268_));
 sky130_fd_sc_hd__and4_1 _10364_ (.A(net1825),
    .B(net43),
    .C(net1713),
    .D(net1926),
    .X(_04269_));
 sky130_fd_sc_hd__inv_2 _10365_ (.A(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__a22o_1 _10366_ (.A1(net731),
    .A2(net869),
    .B1(net1717),
    .B2(net914),
    .X(_04271_));
 sky130_fd_sc_hd__a22o_1 _10367_ (.A1(net43),
    .A2(net1713),
    .B1(net1926),
    .B2(net1825),
    .X(_04272_));
 sky130_fd_sc_hd__or4bb_2 _10368_ (.A(_04251_),
    .B(_04269_),
    .C_N(_04271_),
    .D_N(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a21o_1 _10369_ (.A1(_04270_),
    .A2(_04273_),
    .B1(_04268_),
    .X(_04274_));
 sky130_fd_sc_hd__nand3_1 _10370_ (.A(_04268_),
    .B(_04270_),
    .C(_04273_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand2_1 _10371_ (.A(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__a22o_1 _10372_ (.A1(_04252_),
    .A2(_04271_),
    .B1(_04272_),
    .B2(_04270_),
    .X(_04277_));
 sky130_fd_sc_hd__and4_1 _10373_ (.A(net43),
    .B(net914),
    .C(net1713),
    .D(net1926),
    .X(_04278_));
 sky130_fd_sc_hd__a22o_1 _10374_ (.A1(net914),
    .A2(net1713),
    .B1(net1926),
    .B2(net43),
    .X(_04279_));
 sky130_fd_sc_hd__inv_2 _10375_ (.A(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__and4b_1 _10376_ (.A_N(_04278_),
    .B(_04279_),
    .C(net731),
    .D(net1717),
    .X(_04281_));
 sky130_fd_sc_hd__or2_1 _10377_ (.A(_04278_),
    .B(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__and3_1 _10378_ (.A(_04273_),
    .B(_04277_),
    .C(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__o2bb2a_1 _10379_ (.A1_N(net731),
    .A2_N(net1717),
    .B1(_04278_),
    .B2(_04280_),
    .X(_04284_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(_04281_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__and4_1 _10381_ (.A(net914),
    .B(net731),
    .C(net1713),
    .D(net1926),
    .X(_04286_));
 sky130_fd_sc_hd__and2_2 _10382_ (.A(_04285_),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__a21oi_1 _10383_ (.A1(_04273_),
    .A2(_04277_),
    .B1(_04282_),
    .Y(_04288_));
 sky130_fd_sc_hd__nor2_1 _10384_ (.A(_04283_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__a21oi_2 _10385_ (.A1(_04287_),
    .A2(_04289_),
    .B1(_04283_),
    .Y(_04290_));
 sky130_fd_sc_hd__or2_1 _10386_ (.A(_04276_),
    .B(_04290_),
    .X(_04291_));
 sky130_fd_sc_hd__a21o_1 _10387_ (.A1(_04274_),
    .A2(_04291_),
    .B1(_04267_),
    .X(_04292_));
 sky130_fd_sc_hd__or3_1 _10388_ (.A(_04264_),
    .B(_04266_),
    .C(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__a211o_1 _10389_ (.A1(_04265_),
    .A2(_04293_),
    .B1(_04246_),
    .C1(_04248_),
    .X(_04294_));
 sky130_fd_sc_hd__a211oi_2 _10390_ (.A1(_04247_),
    .A2(_04294_),
    .B1(_04225_),
    .C1(_04226_),
    .Y(_04295_));
 sky130_fd_sc_hd__o21ai_2 _10391_ (.A1(_04225_),
    .A2(_04295_),
    .B1(_04200_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21oi_1 _10392_ (.A1(_04199_),
    .A2(_04296_),
    .B1(_04172_),
    .Y(_04297_));
 sky130_fd_sc_hd__o21a_1 _10393_ (.A1(_04170_),
    .A2(_04297_),
    .B1(_04143_),
    .X(_04298_));
 sky130_fd_sc_hd__o21ba_1 _10394_ (.A1(_04122_),
    .A2(_04142_),
    .B1_N(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__o21a_1 _10395_ (.A1(_04120_),
    .A2(_04299_),
    .B1(_04117_),
    .X(_04300_));
 sky130_fd_sc_hd__xnor2_2 _10396_ (.A(_04091_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21o_1 _10397_ (.A1(_03781_),
    .A2(_04034_),
    .B1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__and2_1 _10398_ (.A(net540),
    .B(net1672),
    .X(_04303_));
 sky130_fd_sc_hd__and3_1 _10399_ (.A(net899),
    .B(net1709),
    .C(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__nand3_1 _10400_ (.A(net899),
    .B(net1709),
    .C(_04303_),
    .Y(_04305_));
 sky130_fd_sc_hd__a22o_1 _10401_ (.A1(net540),
    .A2(net1709),
    .B1(net1672),
    .B2(net1448),
    .X(_04306_));
 sky130_fd_sc_hd__nand4_1 _10402_ (.A(net1448),
    .B(net540),
    .C(net1709),
    .D(net1672),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2_1 _10403_ (.A(_04306_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__a21o_1 _10404_ (.A1(net899),
    .A2(net1709),
    .B1(_04303_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(net540),
    .B(net737),
    .Y(_04310_));
 sky130_fd_sc_hd__and3_1 _10406_ (.A(net1448),
    .B(net1887),
    .C(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__and3_1 _10407_ (.A(_04305_),
    .B(_04309_),
    .C(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__and4_1 _10408_ (.A(net1448),
    .B(net540),
    .C(net1887),
    .D(net2447),
    .X(_04313_));
 sky130_fd_sc_hd__or2_1 _10409_ (.A(_04312_),
    .B(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__nand2b_1 _10410_ (.A_N(_04308_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__xnor2_1 _10411_ (.A(_04308_),
    .B(_04314_),
    .Y(_04316_));
 sky130_fd_sc_hd__xnor2_1 _10412_ (.A(_04304_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__a21oi_1 _10413_ (.A1(_04305_),
    .A2(_04309_),
    .B1(_04311_),
    .Y(_04318_));
 sky130_fd_sc_hd__or2_1 _10414_ (.A(_04312_),
    .B(_04318_),
    .X(_04319_));
 sky130_fd_sc_hd__a22oi_1 _10415_ (.A1(net540),
    .A2(net1887),
    .B1(net737),
    .B2(net1448),
    .Y(_04320_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_04313_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__a22o_1 _10417_ (.A1(net540),
    .A2(net737),
    .B1(net767),
    .B2(net1448),
    .X(_04322_));
 sky130_fd_sc_hd__and4_1 _10418_ (.A(net1448),
    .B(net540),
    .C(net2447),
    .D(net767),
    .X(_04323_));
 sky130_fd_sc_hd__nand4_1 _10419_ (.A(net1448),
    .B(net540),
    .C(net737),
    .D(net767),
    .Y(_04324_));
 sky130_fd_sc_hd__and4_1 _10420_ (.A(net899),
    .B(net1887),
    .C(_04322_),
    .D(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__xnor2_1 _10421_ (.A(_04321_),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__a21oi_1 _10422_ (.A1(net755),
    .A2(net1709),
    .B1(_04323_),
    .Y(_04327_));
 sky130_fd_sc_hd__and3_1 _10423_ (.A(net755),
    .B(net1709),
    .C(_04323_),
    .X(_04328_));
 sky130_fd_sc_hd__or2_1 _10424_ (.A(_04327_),
    .B(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__nand2_1 _10425_ (.A(net899),
    .B(net1672),
    .Y(_04330_));
 sky130_fd_sc_hd__xnor2_1 _10426_ (.A(_04329_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nor2_1 _10427_ (.A(_04326_),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__a21oi_1 _10428_ (.A1(_04321_),
    .A2(_04325_),
    .B1(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__or2_1 _10429_ (.A(_04319_),
    .B(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__xor2_1 _10430_ (.A(_04319_),
    .B(_04333_),
    .X(_04335_));
 sky130_fd_sc_hd__o21bai_1 _10431_ (.A1(_04327_),
    .A2(_04330_),
    .B1_N(_04328_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10432_ (.A(_04335_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__a21o_1 _10433_ (.A1(_04334_),
    .A2(_04337_),
    .B1(_04317_),
    .X(_04338_));
 sky130_fd_sc_hd__nand3_1 _10434_ (.A(_04317_),
    .B(_04334_),
    .C(_04337_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_1 _10435_ (.A(_04338_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__xnor2_1 _10436_ (.A(_04335_),
    .B(_04336_),
    .Y(_04341_));
 sky130_fd_sc_hd__and2_1 _10437_ (.A(_04326_),
    .B(_04331_),
    .X(_04342_));
 sky130_fd_sc_hd__nor2_1 _10438_ (.A(_04332_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__a22oi_1 _10439_ (.A1(net899),
    .A2(net1887),
    .B1(_04322_),
    .B2(_04324_),
    .Y(_04344_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_04325_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__and4_1 _10441_ (.A(net1448),
    .B(net1861),
    .C(net1887),
    .D(net839),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(net755),
    .B(net1887),
    .Y(_04347_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(_04347_),
    .A1(net755),
    .S(_04346_),
    .X(_04348_));
 sky130_fd_sc_hd__a22oi_1 _10444_ (.A1(net899),
    .A2(net737),
    .B1(net767),
    .B2(net540),
    .Y(_04349_));
 sky130_fd_sc_hd__and4_1 _10445_ (.A(net1486),
    .B(net899),
    .C(net737),
    .D(net767),
    .X(_04350_));
 sky130_fd_sc_hd__nor2_1 _10446_ (.A(_04349_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_1 _10447_ (.A(net1448),
    .B(net2189),
    .Y(_04352_));
 sky130_fd_sc_hd__xor2_1 _10448_ (.A(_04351_),
    .B(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__o2bb2a_1 _10449_ (.A1_N(net2487),
    .A2_N(_04346_),
    .B1(_04348_),
    .B2(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__and2b_1 _10450_ (.A_N(_04354_),
    .B(_04345_),
    .X(_04355_));
 sky130_fd_sc_hd__and2b_1 _10451_ (.A_N(_04345_),
    .B(_04354_),
    .X(_04356_));
 sky130_fd_sc_hd__or2_1 _10452_ (.A(_04355_),
    .B(_04356_),
    .X(_04357_));
 sky130_fd_sc_hd__a31o_1 _10453_ (.A1(net1448),
    .A2(net2189),
    .A3(_04351_),
    .B1(_04350_),
    .X(_04358_));
 sky130_fd_sc_hd__and2_1 _10454_ (.A(net1861),
    .B(net1709),
    .X(_04359_));
 sky130_fd_sc_hd__nor2_1 _10455_ (.A(_04358_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__and2_1 _10456_ (.A(_04358_),
    .B(_04359_),
    .X(_04361_));
 sky130_fd_sc_hd__nor2_1 _10457_ (.A(_04360_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(net755),
    .B(net1672),
    .Y(_04363_));
 sky130_fd_sc_hd__xor2_1 _10459_ (.A(_04362_),
    .B(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__nor2_1 _10460_ (.A(_04357_),
    .B(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__o21ai_1 _10461_ (.A1(_04355_),
    .A2(_04365_),
    .B1(_04343_),
    .Y(_04366_));
 sky130_fd_sc_hd__or3_1 _10462_ (.A(_04343_),
    .B(_04355_),
    .C(_04365_),
    .X(_04367_));
 sky130_fd_sc_hd__and2_1 _10463_ (.A(_04366_),
    .B(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o21ba_1 _10464_ (.A1(_04360_),
    .A2(_04363_),
    .B1_N(_04361_),
    .X(_04369_));
 sky130_fd_sc_hd__nand2b_1 _10465_ (.A_N(_04369_),
    .B(_04368_),
    .Y(_04370_));
 sky130_fd_sc_hd__a21o_1 _10466_ (.A1(_04366_),
    .A2(_04370_),
    .B1(_04341_),
    .X(_04371_));
 sky130_fd_sc_hd__nand3_1 _10467_ (.A(_04341_),
    .B(_04366_),
    .C(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _10468_ (.A(_04371_),
    .B(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hd__xnor2_1 _10469_ (.A(_04368_),
    .B(_04369_),
    .Y(_04374_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(_04357_),
    .B(_04364_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand2b_1 _10471_ (.A_N(_04365_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__xor2_1 _10472_ (.A(_04348_),
    .B(_04353_),
    .X(_04377_));
 sky130_fd_sc_hd__a22oi_1 _10473_ (.A1(net1861),
    .A2(net1887),
    .B1(net839),
    .B2(net1448),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_1 _10474_ (.A(_04346_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__and4_1 _10475_ (.A(net1448),
    .B(net540),
    .C(net839),
    .D(net896),
    .X(_04380_));
 sky130_fd_sc_hd__a22o_1 _10476_ (.A1(net540),
    .A2(net839),
    .B1(net896),
    .B2(net1448),
    .X(_04381_));
 sky130_fd_sc_hd__and2b_1 _10477_ (.A_N(_04380_),
    .B(_04381_),
    .X(_04382_));
 sky130_fd_sc_hd__nand2_1 _10478_ (.A(net1686),
    .B(net1887),
    .Y(_04383_));
 sky130_fd_sc_hd__a31o_1 _10479_ (.A1(net1686),
    .A2(net1887),
    .A3(_04381_),
    .B1(_04380_),
    .X(_04384_));
 sky130_fd_sc_hd__and2_1 _10480_ (.A(_04379_),
    .B(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__xnor2_1 _10481_ (.A(_04379_),
    .B(_04384_),
    .Y(_04386_));
 sky130_fd_sc_hd__a22oi_1 _10482_ (.A1(net755),
    .A2(net737),
    .B1(net767),
    .B2(net2493),
    .Y(_04387_));
 sky130_fd_sc_hd__and4_1 _10483_ (.A(net2493),
    .B(net755),
    .C(net737),
    .D(net767),
    .X(_04388_));
 sky130_fd_sc_hd__or2_1 _10484_ (.A(_04387_),
    .B(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__nand2_1 _10485_ (.A(net1486),
    .B(net2189),
    .Y(_04390_));
 sky130_fd_sc_hd__xnor2_1 _10486_ (.A(_04389_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__nor2_1 _10487_ (.A(_04386_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__o21ai_1 _10488_ (.A1(_04385_),
    .A2(_04392_),
    .B1(_04377_),
    .Y(_04393_));
 sky130_fd_sc_hd__or3_1 _10489_ (.A(_04377_),
    .B(_04385_),
    .C(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__and2_1 _10490_ (.A(_04393_),
    .B(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__o21bai_1 _10491_ (.A1(_04387_),
    .A2(_04390_),
    .B1_N(_04388_),
    .Y(_04396_));
 sky130_fd_sc_hd__and2_1 _10492_ (.A(net1686),
    .B(net1709),
    .X(_04397_));
 sky130_fd_sc_hd__nor2_1 _10493_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__and2_1 _10494_ (.A(_04396_),
    .B(_04397_),
    .X(_04399_));
 sky130_fd_sc_hd__nor2_1 _10495_ (.A(_04398_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _10496_ (.A(net1861),
    .B(net1672),
    .Y(_04401_));
 sky130_fd_sc_hd__xnor2_1 _10497_ (.A(_04400_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand2_1 _10498_ (.A(_04395_),
    .B(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__a21oi_1 _10499_ (.A1(_04393_),
    .A2(_04403_),
    .B1(_04376_),
    .Y(_04404_));
 sky130_fd_sc_hd__and3_1 _10500_ (.A(_04376_),
    .B(_04393_),
    .C(_04403_),
    .X(_04405_));
 sky130_fd_sc_hd__or2_1 _10501_ (.A(_04404_),
    .B(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__o21ba_1 _10502_ (.A1(_04398_),
    .A2(_04401_),
    .B1_N(_04399_),
    .X(_04407_));
 sky130_fd_sc_hd__nor2_1 _10503_ (.A(_04406_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__o21ai_1 _10504_ (.A1(_04404_),
    .A2(_04408_),
    .B1(_04374_),
    .Y(_04409_));
 sky130_fd_sc_hd__or3_1 _10505_ (.A(_04374_),
    .B(_04404_),
    .C(_04408_),
    .X(_04410_));
 sky130_fd_sc_hd__and2_1 _10506_ (.A(_04409_),
    .B(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__xnor2_1 _10507_ (.A(_04406_),
    .B(_04407_),
    .Y(_04412_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(_04395_),
    .B(_04402_),
    .X(_04413_));
 sky130_fd_sc_hd__nand2_1 _10509_ (.A(_04403_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__and2_1 _10510_ (.A(_04386_),
    .B(_04391_),
    .X(_04415_));
 sky130_fd_sc_hd__or2_1 _10511_ (.A(_04392_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__xnor2_1 _10512_ (.A(_04382_),
    .B(_04383_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand4_2 _10513_ (.A(net540),
    .B(net899),
    .C(net839),
    .D(net896),
    .Y(_04418_));
 sky130_fd_sc_hd__a22o_1 _10514_ (.A1(net899),
    .A2(net839),
    .B1(net896),
    .B2(net540),
    .X(_04419_));
 sky130_fd_sc_hd__and4_1 _10515_ (.A(net1652),
    .B(net1887),
    .C(_04418_),
    .D(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__a41o_1 _10516_ (.A1(net540),
    .A2(net899),
    .A3(net839),
    .A4(net896),
    .B1(_04420_),
    .X(_04421_));
 sky130_fd_sc_hd__nand2_1 _10517_ (.A(_04417_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__xnor2_1 _10518_ (.A(_04417_),
    .B(_04421_),
    .Y(_04423_));
 sky130_fd_sc_hd__a22oi_1 _10519_ (.A1(net1861),
    .A2(net2447),
    .B1(net767),
    .B2(net755),
    .Y(_04424_));
 sky130_fd_sc_hd__and4_1 _10520_ (.A(net755),
    .B(net1861),
    .C(net2447),
    .D(net2431),
    .X(_04425_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(_04424_),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2_1 _10522_ (.A(net899),
    .B(net2189),
    .Y(_04427_));
 sky130_fd_sc_hd__xor2_1 _10523_ (.A(_04426_),
    .B(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__or2_1 _10524_ (.A(_04423_),
    .B(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__a21o_1 _10525_ (.A1(_04422_),
    .A2(_04429_),
    .B1(_04416_),
    .X(_04430_));
 sky130_fd_sc_hd__nand3_1 _10526_ (.A(_04416_),
    .B(_04422_),
    .C(_04429_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_1 _10527_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__a31o_1 _10528_ (.A1(net899),
    .A2(net2189),
    .A3(_04426_),
    .B1(_04425_),
    .X(_04433_));
 sky130_fd_sc_hd__and2_1 _10529_ (.A(net1652),
    .B(net1709),
    .X(_04434_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(_04433_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__and2_1 _10531_ (.A(_04433_),
    .B(_04434_),
    .X(_04436_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(_04435_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _10533_ (.A(net1686),
    .B(net1672),
    .Y(_04438_));
 sky130_fd_sc_hd__xor2_1 _10534_ (.A(_04437_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__o21a_1 _10535_ (.A1(_04432_),
    .A2(_04439_),
    .B1(_04430_),
    .X(_04440_));
 sky130_fd_sc_hd__xnor2_1 _10536_ (.A(_04414_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__o21ba_1 _10537_ (.A1(_04435_),
    .A2(_04438_),
    .B1_N(_04436_),
    .X(_04442_));
 sky130_fd_sc_hd__or2_1 _10538_ (.A(_04441_),
    .B(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__o21ai_1 _10539_ (.A1(_04414_),
    .A2(_04440_),
    .B1(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__and2b_1 _10540_ (.A_N(_04412_),
    .B(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__xnor2_1 _10541_ (.A(_04412_),
    .B(_04444_),
    .Y(_04446_));
 sky130_fd_sc_hd__xnor2_1 _10542_ (.A(_04441_),
    .B(_04442_),
    .Y(_04447_));
 sky130_fd_sc_hd__xor2_1 _10543_ (.A(_04432_),
    .B(_04439_),
    .X(_04448_));
 sky130_fd_sc_hd__xor2_1 _10544_ (.A(_04423_),
    .B(_04428_),
    .X(_04449_));
 sky130_fd_sc_hd__a22oi_2 _10545_ (.A1(net1652),
    .A2(net1887),
    .B1(_04418_),
    .B2(_04419_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand4_2 _10546_ (.A(net899),
    .B(net755),
    .C(net839),
    .D(net896),
    .Y(_04451_));
 sky130_fd_sc_hd__a22o_1 _10547_ (.A1(net755),
    .A2(net839),
    .B1(net896),
    .B2(net899),
    .X(_04452_));
 sky130_fd_sc_hd__nand4_2 _10548_ (.A(net1574),
    .B(net1887),
    .C(_04451_),
    .D(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__a211oi_2 _10549_ (.A1(_04451_),
    .A2(_04453_),
    .B1(_04420_),
    .C1(_04450_),
    .Y(_04454_));
 sky130_fd_sc_hd__o211a_1 _10550_ (.A1(_04420_),
    .A2(_04450_),
    .B1(_04451_),
    .C1(_04453_),
    .X(_04455_));
 sky130_fd_sc_hd__or2_1 _10551_ (.A(_04454_),
    .B(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__a22oi_1 _10552_ (.A1(net1686),
    .A2(net737),
    .B1(net767),
    .B2(net1861),
    .Y(_04457_));
 sky130_fd_sc_hd__and4_1 _10553_ (.A(net1861),
    .B(net1686),
    .C(net737),
    .D(net767),
    .X(_04458_));
 sky130_fd_sc_hd__nor2_1 _10554_ (.A(_04457_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _10555_ (.A(net755),
    .B(net2189),
    .Y(_04460_));
 sky130_fd_sc_hd__xor2_1 _10556_ (.A(_04459_),
    .B(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__nor2_1 _10557_ (.A(_04456_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21a_1 _10558_ (.A1(_04454_),
    .A2(_04462_),
    .B1(_04449_),
    .X(_04463_));
 sky130_fd_sc_hd__nor3_1 _10559_ (.A(_04449_),
    .B(_04454_),
    .C(_04462_),
    .Y(_04464_));
 sky130_fd_sc_hd__a31o_1 _10560_ (.A1(net755),
    .A2(net2189),
    .A3(_04459_),
    .B1(_04458_),
    .X(_04465_));
 sky130_fd_sc_hd__a21oi_1 _10561_ (.A1(net1574),
    .A2(net1709),
    .B1(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__and3_1 _10562_ (.A(net1574),
    .B(net1709),
    .C(_04465_),
    .X(_04467_));
 sky130_fd_sc_hd__nor2_1 _10563_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_1 _10564_ (.A(net1652),
    .B(net1672),
    .Y(_04469_));
 sky130_fd_sc_hd__xor2_1 _10565_ (.A(_04468_),
    .B(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__or3_1 _10566_ (.A(_04463_),
    .B(_04464_),
    .C(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__and2b_1 _10567_ (.A_N(_04463_),
    .B(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__nand2b_1 _10568_ (.A_N(_04472_),
    .B(_04448_),
    .Y(_04473_));
 sky130_fd_sc_hd__xnor2_1 _10569_ (.A(_04448_),
    .B(_04472_),
    .Y(_04474_));
 sky130_fd_sc_hd__o21ba_1 _10570_ (.A1(_04466_),
    .A2(_04469_),
    .B1_N(_04467_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2b_1 _10571_ (.A_N(_04475_),
    .B(_04474_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21oi_1 _10572_ (.A1(_04473_),
    .A2(_04476_),
    .B1(_04447_),
    .Y(_04477_));
 sky130_fd_sc_hd__and3_1 _10573_ (.A(_04447_),
    .B(_04473_),
    .C(_04476_),
    .X(_04478_));
 sky130_fd_sc_hd__or2_1 _10574_ (.A(_04477_),
    .B(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__xnor2_1 _10575_ (.A(_04474_),
    .B(_04475_),
    .Y(_04480_));
 sky130_fd_sc_hd__o21ai_1 _10576_ (.A1(_04463_),
    .A2(_04464_),
    .B1(_04470_),
    .Y(_04481_));
 sky130_fd_sc_hd__xor2_1 _10577_ (.A(_04456_),
    .B(_04461_),
    .X(_04482_));
 sky130_fd_sc_hd__a22o_1 _10578_ (.A1(net1574),
    .A2(net1887),
    .B1(_04451_),
    .B2(_04452_),
    .X(_04483_));
 sky130_fd_sc_hd__and4_1 _10579_ (.A(net755),
    .B(net1861),
    .C(net839),
    .D(net896),
    .X(_04484_));
 sky130_fd_sc_hd__and3_1 _10580_ (.A(_04453_),
    .B(_04483_),
    .C(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_1 _10581_ (.A1(_04453_),
    .A2(_04483_),
    .B1(_04484_),
    .Y(_04486_));
 sky130_fd_sc_hd__nor2_1 _10582_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a22oi_1 _10583_ (.A1(net1652),
    .A2(net737),
    .B1(net767),
    .B2(net1686),
    .Y(_04488_));
 sky130_fd_sc_hd__and4_1 _10584_ (.A(net1686),
    .B(net1652),
    .C(net737),
    .D(net767),
    .X(_04489_));
 sky130_fd_sc_hd__nor2_1 _10585_ (.A(_04488_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a21oi_1 _10586_ (.A1(net1861),
    .A2(net2189),
    .B1(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__and3_1 _10587_ (.A(net1861),
    .B(net2189),
    .C(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__nor2_1 _10588_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21oi_1 _10589_ (.A1(_04487_),
    .A2(_04493_),
    .B1(_04485_),
    .Y(_04494_));
 sky130_fd_sc_hd__and2b_1 _10590_ (.A_N(_04494_),
    .B(_04482_),
    .X(_04495_));
 sky130_fd_sc_hd__xnor2_1 _10591_ (.A(_04482_),
    .B(_04494_),
    .Y(_04496_));
 sky130_fd_sc_hd__o211a_1 _10592_ (.A1(_04489_),
    .A2(_04492_),
    .B1(net1574),
    .C1(net1672),
    .X(_04497_));
 sky130_fd_sc_hd__a211oi_1 _10593_ (.A1(net1574),
    .A2(net1672),
    .B1(_04489_),
    .C1(_04492_),
    .Y(_04498_));
 sky130_fd_sc_hd__nor2_1 _10594_ (.A(_04497_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__and2_1 _10595_ (.A(_04496_),
    .B(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__o211a_1 _10596_ (.A1(_04495_),
    .A2(_04500_),
    .B1(_04471_),
    .C1(_04481_),
    .X(_04501_));
 sky130_fd_sc_hd__a211o_1 _10597_ (.A1(_04471_),
    .A2(_04481_),
    .B1(_04495_),
    .C1(_04500_),
    .X(_04502_));
 sky130_fd_sc_hd__and2b_1 _10598_ (.A_N(_04501_),
    .B(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__a21oi_1 _10599_ (.A1(_04497_),
    .A2(_04502_),
    .B1(_04501_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2b_1 _10600_ (.A_N(_04504_),
    .B(_04480_),
    .Y(_04505_));
 sky130_fd_sc_hd__xnor2_1 _10601_ (.A(_04480_),
    .B(_04504_),
    .Y(_04506_));
 sky130_fd_sc_hd__xnor2_1 _10602_ (.A(_04497_),
    .B(_04503_),
    .Y(_04507_));
 sky130_fd_sc_hd__nor2_1 _10603_ (.A(_04496_),
    .B(_04499_),
    .Y(_04508_));
 sky130_fd_sc_hd__or2_1 _10604_ (.A(_04500_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_2 _10605_ (.A(_04487_),
    .B(_04493_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand4_2 _10606_ (.A(net1861),
    .B(net1686),
    .C(net839),
    .D(net896),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_1 _10607_ (.A(_04484_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__a22o_1 _10608_ (.A1(net1574),
    .A2(net737),
    .B1(net767),
    .B2(net1652),
    .X(_04513_));
 sky130_fd_sc_hd__and3_1 _10609_ (.A(net1652),
    .B(net1574),
    .C(net767),
    .X(_04514_));
 sky130_fd_sc_hd__a21bo_1 _10610_ (.A1(net737),
    .A2(_04514_),
    .B1_N(_04513_),
    .X(_04515_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(net1686),
    .B(net2189),
    .Y(_04516_));
 sky130_fd_sc_hd__xor2_2 _10612_ (.A(_04515_),
    .B(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__inv_2 _10613_ (.A(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(_04484_),
    .B(_04511_),
    .X(_04519_));
 sky130_fd_sc_hd__a22o_1 _10615_ (.A1(net1861),
    .A2(net839),
    .B1(net896),
    .B2(net755),
    .X(_04520_));
 sky130_fd_sc_hd__or3b_1 _10616_ (.A(_04512_),
    .B(_04519_),
    .C_N(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__o21ba_1 _10617_ (.A1(_04518_),
    .A2(_04521_),
    .B1_N(_04512_),
    .X(_04522_));
 sky130_fd_sc_hd__nor2_1 _10618_ (.A(_04510_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__xor2_2 _10619_ (.A(_04510_),
    .B(_04522_),
    .X(_04524_));
 sky130_fd_sc_hd__a32o_1 _10620_ (.A1(net1686),
    .A2(net2189),
    .A3(_04513_),
    .B1(_04514_),
    .B2(net737),
    .X(_04525_));
 sky130_fd_sc_hd__a21o_1 _10621_ (.A1(_04524_),
    .A2(_04525_),
    .B1(_04523_),
    .X(_04526_));
 sky130_fd_sc_hd__nand2b_1 _10622_ (.A_N(_04509_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__xnor2_1 _10623_ (.A(_04509_),
    .B(_04526_),
    .Y(_04528_));
 sky130_fd_sc_hd__xor2_2 _10624_ (.A(_04524_),
    .B(_04525_),
    .X(_04529_));
 sky130_fd_sc_hd__xor2_1 _10625_ (.A(_04517_),
    .B(_04521_),
    .X(_04530_));
 sky130_fd_sc_hd__nand4_2 _10626_ (.A(net1686),
    .B(net1652),
    .C(net839),
    .D(net896),
    .Y(_04531_));
 sky130_fd_sc_hd__and2b_1 _10627_ (.A_N(_04531_),
    .B(_04511_),
    .X(_04532_));
 sky130_fd_sc_hd__a22o_1 _10628_ (.A1(net1574),
    .A2(net767),
    .B1(net2189),
    .B2(net1652),
    .X(_04533_));
 sky130_fd_sc_hd__nand2_1 _10629_ (.A(net2189),
    .B(_04514_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _10630_ (.A(_04533_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__and2b_1 _10631_ (.A_N(_04511_),
    .B(_04531_),
    .X(_04536_));
 sky130_fd_sc_hd__a22o_1 _10632_ (.A1(net1686),
    .A2(net2425),
    .B1(net896),
    .B2(net1861),
    .X(_04537_));
 sky130_fd_sc_hd__or3b_1 _10633_ (.A(_04532_),
    .B(_04536_),
    .C_N(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__o21bai_1 _10634_ (.A1(_04535_),
    .A2(_04538_),
    .B1_N(_04532_),
    .Y(_04539_));
 sky130_fd_sc_hd__and2b_1 _10635_ (.A_N(_04530_),
    .B(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__xor2_1 _10636_ (.A(_04530_),
    .B(_04539_),
    .X(_04541_));
 sky130_fd_sc_hd__nor2_1 _10637_ (.A(_04534_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__or2_1 _10638_ (.A(_04540_),
    .B(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__and2_1 _10639_ (.A(_04529_),
    .B(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__xnor2_2 _10640_ (.A(_04529_),
    .B(_04543_),
    .Y(_04545_));
 sky130_fd_sc_hd__and2_1 _10641_ (.A(_04534_),
    .B(_04541_),
    .X(_04546_));
 sky130_fd_sc_hd__or2_1 _10642_ (.A(_04542_),
    .B(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__xor2_1 _10643_ (.A(_04535_),
    .B(_04538_),
    .X(_04548_));
 sky130_fd_sc_hd__and4_1 _10644_ (.A(net1652),
    .B(net1574),
    .C(net2425),
    .D(net896),
    .X(_04549_));
 sky130_fd_sc_hd__nand2_1 _10645_ (.A(_04531_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_1 _10646_ (.A(net1574),
    .B(net2189),
    .Y(_04551_));
 sky130_fd_sc_hd__or2_1 _10647_ (.A(_04531_),
    .B(_04549_),
    .X(_04552_));
 sky130_fd_sc_hd__a22o_1 _10648_ (.A1(net1652),
    .A2(net2427),
    .B1(net2007),
    .B2(net1686),
    .X(_04553_));
 sky130_fd_sc_hd__nand3_2 _10649_ (.A(_04550_),
    .B(_04552_),
    .C(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__o21ai_1 _10650_ (.A1(_04551_),
    .A2(_04554_),
    .B1(_04550_),
    .Y(_04555_));
 sky130_fd_sc_hd__and2_1 _10651_ (.A(_04548_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__and2b_1 _10652_ (.A_N(_04547_),
    .B(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__and2b_1 _10653_ (.A_N(_04545_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__o21ai_1 _10654_ (.A1(_04544_),
    .A2(_04558_),
    .B1(_04528_),
    .Y(_04559_));
 sky130_fd_sc_hd__a21oi_1 _10655_ (.A1(_04527_),
    .A2(_04559_),
    .B1(_04507_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _10656_ (.A(_04506_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__a21oi_1 _10657_ (.A1(_04505_),
    .A2(_04561_),
    .B1(_04479_),
    .Y(_04562_));
 sky130_fd_sc_hd__o21a_1 _10658_ (.A1(_04477_),
    .A2(_04562_),
    .B1(_04446_),
    .X(_04563_));
 sky130_fd_sc_hd__o21ai_1 _10659_ (.A1(_04445_),
    .A2(_04563_),
    .B1(_04411_),
    .Y(_04564_));
 sky130_fd_sc_hd__a21o_1 _10660_ (.A1(_04409_),
    .A2(_04564_),
    .B1(_04373_),
    .X(_04565_));
 sky130_fd_sc_hd__a21o_1 _10661_ (.A1(_04371_),
    .A2(_04565_),
    .B1(_04340_),
    .X(_04566_));
 sky130_fd_sc_hd__nand3_1 _10662_ (.A(_04340_),
    .B(_04371_),
    .C(_04565_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand2_2 _10663_ (.A(_04566_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand3_1 _10664_ (.A(_03781_),
    .B(_04034_),
    .C(_04301_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand2_1 _10665_ (.A(_04302_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__o21ai_1 _10666_ (.A1(_04568_),
    .A2(_04570_),
    .B1(_04302_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21bo_1 _10667_ (.A1(_04304_),
    .A2(_04316_),
    .B1_N(_04315_),
    .X(_04572_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(net1448),
    .B(net1709),
    .Y(_04573_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(_04303_),
    .B(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__xnor2_1 _10670_ (.A(_04572_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21oi_1 _10671_ (.A1(_04338_),
    .A2(_04566_),
    .B1(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__and3_1 _10672_ (.A(_04338_),
    .B(_04566_),
    .C(_04575_),
    .X(_04577_));
 sky130_fd_sc_hd__nor2_2 _10673_ (.A(_04576_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__a22oi_1 _10674_ (.A1(net421),
    .A2(net1898),
    .B1(net462),
    .B2(net1381),
    .Y(_04579_));
 sky130_fd_sc_hd__and4_1 _10675_ (.A(net1381),
    .B(net421),
    .C(net1898),
    .D(net462),
    .X(_04580_));
 sky130_fd_sc_hd__nor2_1 _10676_ (.A(_04579_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__a32o_1 _10677_ (.A1(net1381),
    .A2(net1747),
    .A3(_03277_),
    .B1(_03278_),
    .B2(net421),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_1 _10678_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__or2_1 _10679_ (.A(_04581_),
    .B(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__nand2_2 _10680_ (.A(_04583_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_03286_),
    .B(_03301_),
    .Y(_04586_));
 sky130_fd_sc_hd__xnor2_2 _10682_ (.A(_04585_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2b_1 _10683_ (.A_N(_03319_),
    .B(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__xnor2_2 _10684_ (.A(_03319_),
    .B(_04587_),
    .Y(_04589_));
 sky130_fd_sc_hd__o21ai_4 _10685_ (.A1(_03344_),
    .A2(_03525_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__or3_4 _10686_ (.A(_03344_),
    .B(_03525_),
    .C(_04589_),
    .X(_04591_));
 sky130_fd_sc_hd__a22oi_1 _10687_ (.A1(net51),
    .A2(net1991),
    .B1(net686),
    .B2(net1425),
    .Y(_04592_));
 sky130_fd_sc_hd__and4_1 _10688_ (.A(net1425),
    .B(net51),
    .C(net1991),
    .D(net686),
    .X(_04593_));
 sky130_fd_sc_hd__nor2_1 _10689_ (.A(_04592_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__a32o_1 _10690_ (.A1(net1425),
    .A2(net1845),
    .A3(_03529_),
    .B1(_03530_),
    .B2(net51),
    .X(_04595_));
 sky130_fd_sc_hd__nand2_1 _10691_ (.A(_04594_),
    .B(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__or2_1 _10692_ (.A(_04594_),
    .B(_04595_),
    .X(_04597_));
 sky130_fd_sc_hd__nand2_2 _10693_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _10694_ (.A(_03538_),
    .B(_03553_),
    .Y(_04599_));
 sky130_fd_sc_hd__xnor2_2 _10695_ (.A(_04598_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2b_1 _10696_ (.A_N(_03571_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__xnor2_2 _10697_ (.A(_03571_),
    .B(_04600_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_4 _10698_ (.A1(_03596_),
    .A2(_03778_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__or3_2 _10699_ (.A(_03596_),
    .B(_03778_),
    .C(_04602_),
    .X(_04604_));
 sky130_fd_sc_hd__nand4_1 _10700_ (.A(_04590_),
    .B(_04591_),
    .C(_04603_),
    .D(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a22oi_1 _10701_ (.A1(net440),
    .A2(net1857),
    .B1(net675),
    .B2(net1393),
    .Y(_04606_));
 sky130_fd_sc_hd__and4_1 _10702_ (.A(net1393),
    .B(net440),
    .C(net1857),
    .D(net675),
    .X(_04607_));
 sky130_fd_sc_hd__nor2_1 _10703_ (.A(_04606_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__a32o_1 _10704_ (.A1(net1393),
    .A2(net1870),
    .A3(_03783_),
    .B1(_03784_),
    .B2(net932),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_1 _10705_ (.A(_04608_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__or2_1 _10706_ (.A(_04608_),
    .B(_04609_),
    .X(_04611_));
 sky130_fd_sc_hd__nand2_1 _10707_ (.A(_04610_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__nand2_1 _10708_ (.A(_03793_),
    .B(_03807_),
    .Y(_04613_));
 sky130_fd_sc_hd__xnor2_1 _10709_ (.A(_04612_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2b_1 _10710_ (.A_N(_03826_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__xnor2_1 _10711_ (.A(_03826_),
    .B(_04614_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21ai_2 _10712_ (.A1(_03851_),
    .A2(_04030_),
    .B1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__or3_1 _10713_ (.A(_03851_),
    .B(_04030_),
    .C(_04616_),
    .X(_04618_));
 sky130_fd_sc_hd__a22o_1 _10714_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04603_),
    .B2(_04604_),
    .X(_04619_));
 sky130_fd_sc_hd__and4_1 _10715_ (.A(_04605_),
    .B(_04617_),
    .C(_04618_),
    .D(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__a41o_1 _10716_ (.A1(_04590_),
    .A2(_04591_),
    .A3(_04603_),
    .A4(_04604_),
    .B1(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__and3_1 _10717_ (.A(net1429),
    .B(net1930),
    .C(_04035_),
    .X(_04622_));
 sky130_fd_sc_hd__o21ai_2 _10718_ (.A1(_04046_),
    .A2(_04085_),
    .B1(_04083_),
    .Y(_04623_));
 sky130_fd_sc_hd__xor2_2 _10719_ (.A(_04622_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__nor2_1 _10720_ (.A(_04060_),
    .B(_04085_),
    .Y(_04625_));
 sky130_fd_sc_hd__xnor2_2 _10721_ (.A(_04624_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__o21a_1 _10722_ (.A1(_04091_),
    .A2(_04300_),
    .B1(_04088_),
    .X(_04627_));
 sky130_fd_sc_hd__nor2_1 _10723_ (.A(_04626_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__xnor2_2 _10724_ (.A(_04626_),
    .B(_04627_),
    .Y(_04629_));
 sky130_fd_sc_hd__and2b_1 _10725_ (.A_N(_04629_),
    .B(_04621_),
    .X(_04630_));
 sky130_fd_sc_hd__xnor2_2 _10726_ (.A(_04621_),
    .B(_04629_),
    .Y(_04631_));
 sky130_fd_sc_hd__xnor2_2 _10727_ (.A(_04578_),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__and3_1 _10728_ (.A(net1393),
    .B(net1857),
    .C(_03782_),
    .X(_04633_));
 sky130_fd_sc_hd__o21ai_1 _10729_ (.A1(_03793_),
    .A2(_04612_),
    .B1(_04610_),
    .Y(_04634_));
 sky130_fd_sc_hd__xor2_1 _10730_ (.A(_04633_),
    .B(_04634_),
    .X(_04635_));
 sky130_fd_sc_hd__nor2_1 _10731_ (.A(_03807_),
    .B(_04612_),
    .Y(_04636_));
 sky130_fd_sc_hd__xnor2_1 _10732_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__a21oi_2 _10733_ (.A1(_04615_),
    .A2(_04617_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__and3_1 _10734_ (.A(_04615_),
    .B(_04617_),
    .C(_04637_),
    .X(_04639_));
 sky130_fd_sc_hd__and3_1 _10735_ (.A(net1381),
    .B(net1898),
    .C(_03276_),
    .X(_04640_));
 sky130_fd_sc_hd__o21ai_2 _10736_ (.A1(_03286_),
    .A2(_04585_),
    .B1(_04583_),
    .Y(_04641_));
 sky130_fd_sc_hd__xor2_1 _10737_ (.A(_04640_),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__nor2_1 _10738_ (.A(_03301_),
    .B(_04585_),
    .Y(_04643_));
 sky130_fd_sc_hd__xnor2_1 _10739_ (.A(_04642_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__a21o_2 _10740_ (.A1(_04588_),
    .A2(_04590_),
    .B1(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__nand3_2 _10741_ (.A(_04588_),
    .B(_04590_),
    .C(_04644_),
    .Y(_04646_));
 sky130_fd_sc_hd__and3_1 _10742_ (.A(net1425),
    .B(net1991),
    .C(_03528_),
    .X(_04647_));
 sky130_fd_sc_hd__o21ai_1 _10743_ (.A1(_03538_),
    .A2(_04598_),
    .B1(_04596_),
    .Y(_04648_));
 sky130_fd_sc_hd__xor2_1 _10744_ (.A(_04647_),
    .B(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__nor2_1 _10745_ (.A(_03553_),
    .B(_04598_),
    .Y(_04650_));
 sky130_fd_sc_hd__xnor2_1 _10746_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__a21o_1 _10747_ (.A1(_04601_),
    .A2(_04603_),
    .B1(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__nand3_2 _10748_ (.A(_04601_),
    .B(_04603_),
    .C(_04651_),
    .Y(_04653_));
 sky130_fd_sc_hd__and4_2 _10749_ (.A(_04645_),
    .B(_04646_),
    .C(_04652_),
    .D(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__a22oi_4 _10750_ (.A1(_04645_),
    .A2(_04646_),
    .B1(_04652_),
    .B2(_04653_),
    .Y(_04655_));
 sky130_fd_sc_hd__or4_2 _10751_ (.A(_04638_),
    .B(_04639_),
    .C(_04654_),
    .D(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__o22ai_2 _10752_ (.A1(_04638_),
    .A2(_04639_),
    .B1(_04654_),
    .B2(_04655_),
    .Y(_04657_));
 sky130_fd_sc_hd__and4_1 _10753_ (.A(net557),
    .B(net797),
    .C(net2037),
    .D(net132),
    .X(_04658_));
 sky130_fd_sc_hd__nand4_1 _10754_ (.A(net3664),
    .B(net797),
    .C(net2037),
    .D(net3050),
    .Y(_04659_));
 sky130_fd_sc_hd__nand4_2 _10755_ (.A(net797),
    .B(net953),
    .C(net2037),
    .D(net132),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_1 _10756_ (.A(_04658_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_1 _10757_ (.A(net1438),
    .B(net1987),
    .Y(_04662_));
 sky130_fd_sc_hd__and2_1 _10758_ (.A(_04658_),
    .B(_04660_),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_1 _10759_ (.A1(net797),
    .A2(net2037),
    .B1(net132),
    .B2(net557),
    .X(_04664_));
 sky130_fd_sc_hd__or3b_1 _10760_ (.A(_04661_),
    .B(_04663_),
    .C_N(_04664_),
    .X(_04665_));
 sky130_fd_sc_hd__o21bai_1 _10761_ (.A1(_04662_),
    .A2(_04665_),
    .B1_N(_04661_),
    .Y(_04666_));
 sky130_fd_sc_hd__and4_1 _10762_ (.A(net1438),
    .B(net557),
    .C(net2037),
    .D(net3050),
    .X(_04667_));
 sky130_fd_sc_hd__a22o_1 _10763_ (.A1(net3664),
    .A2(net2037),
    .B1(net132),
    .B2(net1438),
    .X(_04668_));
 sky130_fd_sc_hd__and2_1 _10764_ (.A(_04659_),
    .B(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(_04669_),
    .A1(_04658_),
    .S(_04667_),
    .X(_04670_));
 sky130_fd_sc_hd__nand2_1 _10766_ (.A(_04666_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__nand2_1 _10767_ (.A(net1438),
    .B(net2037),
    .Y(_04672_));
 sky130_fd_sc_hd__a32o_1 _10768_ (.A1(net1438),
    .A2(net557),
    .A3(net3050),
    .B1(net3665),
    .B2(_04672_),
    .X(_04673_));
 sky130_fd_sc_hd__nor2_1 _10769_ (.A(_04671_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__and2_1 _10770_ (.A(_04671_),
    .B(_04673_),
    .X(_04675_));
 sky130_fd_sc_hd__nor2_1 _10771_ (.A(_04674_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__or2_1 _10772_ (.A(_04666_),
    .B(_04670_),
    .X(_04677_));
 sky130_fd_sc_hd__and2_1 _10773_ (.A(_04671_),
    .B(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__xor2_1 _10774_ (.A(_04662_),
    .B(_04665_),
    .X(_04679_));
 sky130_fd_sc_hd__a22o_1 _10775_ (.A1(net953),
    .A2(net2037),
    .B1(net132),
    .B2(net797),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_1 _10776_ (.A1(net953),
    .A2(net132),
    .B1(net992),
    .B2(net1438),
    .X(_04681_));
 sky130_fd_sc_hd__and4_1 _10777_ (.A(net1438),
    .B(net953),
    .C(net132),
    .D(net992),
    .X(_04682_));
 sky130_fd_sc_hd__nand4_1 _10778_ (.A(net1438),
    .B(net2251),
    .C(net132),
    .D(net992),
    .Y(_04683_));
 sky130_fd_sc_hd__and4_1 _10779_ (.A(net69),
    .B(net2037),
    .C(_04681_),
    .D(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__and3_1 _10780_ (.A(_04660_),
    .B(_04680_),
    .C(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__a21oi_1 _10781_ (.A1(_04660_),
    .A2(_04680_),
    .B1(_04684_),
    .Y(_04686_));
 sky130_fd_sc_hd__or2_1 _10782_ (.A(_04685_),
    .B(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_1 _10783_ (.A1(net557),
    .A2(net1987),
    .B1(_04682_),
    .Y(_04688_));
 sky130_fd_sc_hd__and3_1 _10784_ (.A(net557),
    .B(net1987),
    .C(_04682_),
    .X(_04689_));
 sky130_fd_sc_hd__or2_1 _10785_ (.A(_04688_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__nand2_1 _10786_ (.A(net1438),
    .B(net1983),
    .Y(_04691_));
 sky130_fd_sc_hd__xor2_1 _10787_ (.A(_04690_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__and2b_1 _10788_ (.A_N(_04687_),
    .B(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__o21a_1 _10789_ (.A1(_04685_),
    .A2(_04693_),
    .B1(_04679_),
    .X(_04694_));
 sky130_fd_sc_hd__nor3_1 _10790_ (.A(_04679_),
    .B(_04685_),
    .C(_04693_),
    .Y(_04695_));
 sky130_fd_sc_hd__nor2_1 _10791_ (.A(_04694_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__o21ba_1 _10792_ (.A1(_04688_),
    .A2(_04691_),
    .B1_N(_04689_),
    .X(_04697_));
 sky130_fd_sc_hd__and2b_1 _10793_ (.A_N(_04697_),
    .B(_04696_),
    .X(_04698_));
 sky130_fd_sc_hd__o21a_1 _10794_ (.A1(_04694_),
    .A2(_04698_),
    .B1(_04678_),
    .X(_04699_));
 sky130_fd_sc_hd__nor3_1 _10795_ (.A(_04678_),
    .B(_04694_),
    .C(_04698_),
    .Y(_04700_));
 sky130_fd_sc_hd__nor2_1 _10796_ (.A(_04699_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__xnor2_1 _10797_ (.A(_04696_),
    .B(_04697_),
    .Y(_04702_));
 sky130_fd_sc_hd__xor2_1 _10798_ (.A(_04687_),
    .B(_04692_),
    .X(_04703_));
 sky130_fd_sc_hd__a22oi_2 _10799_ (.A1(net69),
    .A2(net2037),
    .B1(_04681_),
    .B2(_04683_),
    .Y(_04704_));
 sky130_fd_sc_hd__nor2_1 _10800_ (.A(_04684_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__and4_1 _10801_ (.A(net1438),
    .B(net1934),
    .C(net2037),
    .D(net1007),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _10802_ (.A(net917),
    .B(net2037),
    .Y(_04707_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(_04707_),
    .A1(net917),
    .S(_04706_),
    .X(_04708_));
 sky130_fd_sc_hd__a22oi_1 _10804_ (.A1(net69),
    .A2(net132),
    .B1(net1970),
    .B2(net1438),
    .Y(_04709_));
 sky130_fd_sc_hd__and4_1 _10805_ (.A(net1438),
    .B(net69),
    .C(net132),
    .D(net1970),
    .X(_04710_));
 sky130_fd_sc_hd__nor2_1 _10806_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _10807_ (.A(net557),
    .B(net992),
    .Y(_04712_));
 sky130_fd_sc_hd__xor2_1 _10808_ (.A(_04711_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__o2bb2a_1 _10809_ (.A1_N(net917),
    .A2_N(_04706_),
    .B1(_04708_),
    .B2(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__or3_1 _10810_ (.A(_04684_),
    .B(_04704_),
    .C(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__xnor2_1 _10811_ (.A(_04705_),
    .B(_04714_),
    .Y(_04716_));
 sky130_fd_sc_hd__a31o_1 _10812_ (.A1(net557),
    .A2(net992),
    .A3(_04711_),
    .B1(_04710_),
    .X(_04717_));
 sky130_fd_sc_hd__and2_1 _10813_ (.A(net3737),
    .B(net1987),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _10814_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__and2_1 _10815_ (.A(_04717_),
    .B(_04718_),
    .X(_04720_));
 sky130_fd_sc_hd__nor2_1 _10816_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _10817_ (.A(net557),
    .B(net1983),
    .Y(_04722_));
 sky130_fd_sc_hd__xnor2_1 _10818_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(_04716_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__a21oi_2 _10820_ (.A1(_04715_),
    .A2(_04724_),
    .B1(_04703_),
    .Y(_04725_));
 sky130_fd_sc_hd__and3_1 _10821_ (.A(_04703_),
    .B(_04715_),
    .C(_04724_),
    .X(_04726_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__o21ba_1 _10823_ (.A1(_04719_),
    .A2(_04722_),
    .B1_N(_04720_),
    .X(_04728_));
 sky130_fd_sc_hd__and2b_1 _10824_ (.A_N(_04728_),
    .B(_04727_),
    .X(_04729_));
 sky130_fd_sc_hd__o21a_1 _10825_ (.A1(_04725_),
    .A2(_04729_),
    .B1(_04702_),
    .X(_04730_));
 sky130_fd_sc_hd__nor3_1 _10826_ (.A(_04702_),
    .B(_04725_),
    .C(_04729_),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _10827_ (.A(_04730_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__xnor2_1 _10828_ (.A(_04727_),
    .B(_04728_),
    .Y(_04733_));
 sky130_fd_sc_hd__or2_1 _10829_ (.A(_04716_),
    .B(_04723_),
    .X(_04734_));
 sky130_fd_sc_hd__nand2_1 _10830_ (.A(_04724_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__xor2_1 _10831_ (.A(_04708_),
    .B(_04713_),
    .X(_04736_));
 sky130_fd_sc_hd__a22oi_1 _10832_ (.A1(net1934),
    .A2(net2037),
    .B1(net1007),
    .B2(net1438),
    .Y(_04737_));
 sky130_fd_sc_hd__or2_1 _10833_ (.A(_04706_),
    .B(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__nand4_1 _10834_ (.A(net1438),
    .B(net557),
    .C(net1007),
    .D(net1010),
    .Y(_04739_));
 sky130_fd_sc_hd__and2_1 _10835_ (.A(net1615),
    .B(net2037),
    .X(_04740_));
 sky130_fd_sc_hd__a22o_1 _10836_ (.A1(net557),
    .A2(net1007),
    .B1(net1010),
    .B2(net1438),
    .X(_04741_));
 sky130_fd_sc_hd__nand3_1 _10837_ (.A(_04739_),
    .B(_04740_),
    .C(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21bo_1 _10838_ (.A1(_04740_),
    .A2(_04741_),
    .B1_N(_04739_),
    .X(_04743_));
 sky130_fd_sc_hd__and2b_1 _10839_ (.A_N(_04738_),
    .B(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__and4_1 _10840_ (.A(net557),
    .B(net917),
    .C(net132),
    .D(net1970),
    .X(_04745_));
 sky130_fd_sc_hd__a22oi_1 _10841_ (.A1(net916),
    .A2(net132),
    .B1(net1970),
    .B2(net557),
    .Y(_04746_));
 sky130_fd_sc_hd__and4bb_1 _10842_ (.A_N(_04745_),
    .B_N(_04746_),
    .C(net797),
    .D(net992),
    .X(_04747_));
 sky130_fd_sc_hd__o2bb2a_1 _10843_ (.A1_N(net797),
    .A2_N(net992),
    .B1(_04745_),
    .B2(_04746_),
    .X(_04748_));
 sky130_fd_sc_hd__nor2_1 _10844_ (.A(_04747_),
    .B(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__xnor2_1 _10845_ (.A(_04738_),
    .B(_04743_),
    .Y(_04750_));
 sky130_fd_sc_hd__and2_1 _10846_ (.A(_04749_),
    .B(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__o21ai_1 _10847_ (.A1(_04744_),
    .A2(_04751_),
    .B1(_04736_),
    .Y(_04752_));
 sky130_fd_sc_hd__or2_2 _10848_ (.A(_04745_),
    .B(_04747_),
    .X(_04753_));
 sky130_fd_sc_hd__nand2_1 _10849_ (.A(net2251),
    .B(net1987),
    .Y(_04754_));
 sky130_fd_sc_hd__xnor2_1 _10850_ (.A(_04753_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__and3_1 _10851_ (.A(net797),
    .B(net1983),
    .C(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__a21oi_1 _10852_ (.A1(net797),
    .A2(net1983),
    .B1(_04755_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor2_1 _10853_ (.A(_04756_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__or3_1 _10854_ (.A(_04736_),
    .B(_04744_),
    .C(_04751_),
    .X(_04759_));
 sky130_fd_sc_hd__and2_1 _10855_ (.A(_04752_),
    .B(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__a21bo_1 _10856_ (.A1(_04758_),
    .A2(_04759_),
    .B1_N(_04752_),
    .X(_04761_));
 sky130_fd_sc_hd__and3_1 _10857_ (.A(_04724_),
    .B(_04734_),
    .C(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__a31oi_4 _10858_ (.A1(net2251),
    .A2(net1987),
    .A3(_04753_),
    .B1(_04756_),
    .Y(_04763_));
 sky130_fd_sc_hd__xor2_2 _10859_ (.A(_04735_),
    .B(_04761_),
    .X(_04764_));
 sky130_fd_sc_hd__nor2_1 _10860_ (.A(_04763_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__or3_2 _10861_ (.A(_04733_),
    .B(_04762_),
    .C(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__o21a_1 _10862_ (.A1(_04762_),
    .A2(_04765_),
    .B1(_04733_),
    .X(_04767_));
 sky130_fd_sc_hd__o21ai_1 _10863_ (.A1(_04762_),
    .A2(_04765_),
    .B1(_04733_),
    .Y(_04768_));
 sky130_fd_sc_hd__xnor2_2 _10864_ (.A(_04763_),
    .B(_04764_),
    .Y(_04769_));
 sky130_fd_sc_hd__xor2_2 _10865_ (.A(_04758_),
    .B(_04760_),
    .X(_04770_));
 sky130_fd_sc_hd__xnor2_1 _10866_ (.A(_04749_),
    .B(_04750_),
    .Y(_04771_));
 sky130_fd_sc_hd__a21o_1 _10867_ (.A1(_04739_),
    .A2(_04741_),
    .B1(_04740_),
    .X(_04772_));
 sky130_fd_sc_hd__and4_1 _10868_ (.A(net557),
    .B(net797),
    .C(net1007),
    .D(net1010),
    .X(_04773_));
 sky130_fd_sc_hd__nand3_1 _10869_ (.A(_04742_),
    .B(_04772_),
    .C(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _10870_ (.A(net953),
    .B(net992),
    .Y(_04775_));
 sky130_fd_sc_hd__a22oi_1 _10871_ (.A1(net1934),
    .A2(net132),
    .B1(net1970),
    .B2(net797),
    .Y(_04776_));
 sky130_fd_sc_hd__and4_1 _10872_ (.A(net797),
    .B(net1934),
    .C(net132),
    .D(net1970),
    .X(_04777_));
 sky130_fd_sc_hd__nor2_1 _10873_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _10874_ (.A(_04775_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__a21o_1 _10875_ (.A1(_04742_),
    .A2(_04772_),
    .B1(_04773_),
    .X(_04780_));
 sky130_fd_sc_hd__nand3_1 _10876_ (.A(_04774_),
    .B(_04779_),
    .C(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__a21bo_1 _10877_ (.A1(_04779_),
    .A2(_04780_),
    .B1_N(_04774_),
    .X(_04782_));
 sky130_fd_sc_hd__and2b_1 _10878_ (.A_N(_04771_),
    .B(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__a31o_1 _10879_ (.A1(net953),
    .A2(net992),
    .A3(_04778_),
    .B1(_04777_),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_1 _10880_ (.A(net1357),
    .B(net1987),
    .Y(_04785_));
 sky130_fd_sc_hd__and3_1 _10881_ (.A(net1357),
    .B(net1987),
    .C(_04784_),
    .X(_04786_));
 sky130_fd_sc_hd__xnor2_1 _10882_ (.A(_04784_),
    .B(_04785_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_1 _10883_ (.A(net953),
    .B(net1983),
    .Y(_04788_));
 sky130_fd_sc_hd__xor2_1 _10884_ (.A(_04787_),
    .B(_04788_),
    .X(_04789_));
 sky130_fd_sc_hd__xor2_1 _10885_ (.A(_04771_),
    .B(_04782_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _10886_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_1 _10887_ (.A(_04783_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__and2b_1 _10888_ (.A_N(_04792_),
    .B(_04770_),
    .X(_04793_));
 sky130_fd_sc_hd__a31o_1 _10889_ (.A1(net953),
    .A2(net1983),
    .A3(_04787_),
    .B1(_04786_),
    .X(_04794_));
 sky130_fd_sc_hd__xnor2_2 _10890_ (.A(_04770_),
    .B(_04792_),
    .Y(_04795_));
 sky130_fd_sc_hd__a21oi_2 _10891_ (.A1(_04794_),
    .A2(_04795_),
    .B1(_04793_),
    .Y(_04796_));
 sky130_fd_sc_hd__nor2_1 _10892_ (.A(_04769_),
    .B(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__xor2_2 _10893_ (.A(_04769_),
    .B(_04796_),
    .X(_04798_));
 sky130_fd_sc_hd__xnor2_2 _10894_ (.A(_04794_),
    .B(_04795_),
    .Y(_04799_));
 sky130_fd_sc_hd__and2_1 _10895_ (.A(_04789_),
    .B(_04790_),
    .X(_04800_));
 sky130_fd_sc_hd__or2_1 _10896_ (.A(_04791_),
    .B(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a21o_1 _10897_ (.A1(_04774_),
    .A2(_04780_),
    .B1(_04779_),
    .X(_04802_));
 sky130_fd_sc_hd__and4_2 _10898_ (.A(net797),
    .B(net953),
    .C(net1007),
    .D(net1010),
    .X(_04803_));
 sky130_fd_sc_hd__inv_2 _10899_ (.A(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__and4_1 _10900_ (.A(net953),
    .B(net1615),
    .C(net132),
    .D(net1970),
    .X(_04805_));
 sky130_fd_sc_hd__a22oi_1 _10901_ (.A1(net1615),
    .A2(net132),
    .B1(net1970),
    .B2(net953),
    .Y(_04806_));
 sky130_fd_sc_hd__and4bb_1 _10902_ (.A_N(_04805_),
    .B_N(_04806_),
    .C(net69),
    .D(net991),
    .X(_04807_));
 sky130_fd_sc_hd__o2bb2a_1 _10903_ (.A1_N(net69),
    .A2_N(net991),
    .B1(_04805_),
    .B2(_04806_),
    .X(_04808_));
 sky130_fd_sc_hd__a22o_1 _10904_ (.A1(net797),
    .A2(net1006),
    .B1(net1010),
    .B2(net557),
    .X(_04809_));
 sky130_fd_sc_hd__xnor2_1 _10905_ (.A(_04773_),
    .B(_04803_),
    .Y(_04810_));
 sky130_fd_sc_hd__or4bb_1 _10906_ (.A(_04807_),
    .B(_04808_),
    .C_N(_04809_),
    .D_N(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__o21ai_1 _10907_ (.A1(_04773_),
    .A2(_04804_),
    .B1(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand3_1 _10908_ (.A(_04781_),
    .B(_04802_),
    .C(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__o211a_1 _10909_ (.A1(_04805_),
    .A2(_04807_),
    .B1(net916),
    .C1(net1987),
    .X(_04814_));
 sky130_fd_sc_hd__a211oi_1 _10910_ (.A1(net916),
    .A2(net1987),
    .B1(_04805_),
    .C1(_04807_),
    .Y(_04815_));
 sky130_fd_sc_hd__nor2_1 _10911_ (.A(net3211),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _10912_ (.A(net69),
    .B(net1983),
    .Y(_04817_));
 sky130_fd_sc_hd__xnor2_1 _10913_ (.A(_04816_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__a21o_1 _10914_ (.A1(_04781_),
    .A2(_04802_),
    .B1(_04812_),
    .X(_04819_));
 sky130_fd_sc_hd__nand3_1 _10915_ (.A(_04813_),
    .B(_04818_),
    .C(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__and2_1 _10916_ (.A(_04813_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__or2_1 _10917_ (.A(_04801_),
    .B(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__a31o_1 _10918_ (.A1(net69),
    .A2(net1983),
    .A3(_04816_),
    .B1(net3211),
    .X(_04823_));
 sky130_fd_sc_hd__xor2_1 _10919_ (.A(_04801_),
    .B(_04821_),
    .X(_04824_));
 sky130_fd_sc_hd__nand2_1 _10920_ (.A(net3212),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__and3_1 _10921_ (.A(_04799_),
    .B(_04822_),
    .C(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__nand3_2 _10922_ (.A(_04799_),
    .B(_04822_),
    .C(_04825_),
    .Y(_04827_));
 sky130_fd_sc_hd__a21oi_1 _10923_ (.A1(_04822_),
    .A2(_04825_),
    .B1(_04799_),
    .Y(_04828_));
 sky130_fd_sc_hd__xnor2_1 _10924_ (.A(net3212),
    .B(_04824_),
    .Y(_04829_));
 sky130_fd_sc_hd__a21o_1 _10925_ (.A1(_04813_),
    .A2(_04819_),
    .B1(_04818_),
    .X(_04830_));
 sky130_fd_sc_hd__a2bb2o_1 _10926_ (.A1_N(_04807_),
    .A2_N(_04808_),
    .B1(_04809_),
    .B2(_04810_),
    .X(_04831_));
 sky130_fd_sc_hd__and4_1 _10927_ (.A(net953),
    .B(net69),
    .C(net1007),
    .D(net1010),
    .X(_04832_));
 sky130_fd_sc_hd__nand4_2 _10928_ (.A(net953),
    .B(net69),
    .C(net1006),
    .D(net1010),
    .Y(_04833_));
 sky130_fd_sc_hd__nor2_1 _10929_ (.A(_04803_),
    .B(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(_04803_),
    .B(_04833_),
    .X(_04835_));
 sky130_fd_sc_hd__a22oi_1 _10931_ (.A1(net917),
    .A2(net992),
    .B1(net1970),
    .B2(net69),
    .Y(_04836_));
 sky130_fd_sc_hd__and4_1 _10932_ (.A(net69),
    .B(net917),
    .C(net992),
    .D(net1970),
    .X(_04837_));
 sky130_fd_sc_hd__nor2_1 _10933_ (.A(_04836_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _10934_ (.A(_04803_),
    .B(_04833_),
    .Y(_04839_));
 sky130_fd_sc_hd__a22o_1 _10935_ (.A1(net953),
    .A2(net1006),
    .B1(net1009),
    .B2(net797),
    .X(_04840_));
 sky130_fd_sc_hd__nand4_1 _10936_ (.A(_04835_),
    .B(_04838_),
    .C(_04839_),
    .D(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__a31o_1 _10937_ (.A1(_04838_),
    .A2(_04839_),
    .A3(_04840_),
    .B1(_04834_),
    .X(_04842_));
 sky130_fd_sc_hd__nand3_1 _10938_ (.A(_04811_),
    .B(_04831_),
    .C(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__a21oi_1 _10939_ (.A1(net1934),
    .A2(net1987),
    .B1(_04837_),
    .Y(_04844_));
 sky130_fd_sc_hd__and3_1 _10940_ (.A(net1934),
    .B(net1987),
    .C(_04837_),
    .X(_04845_));
 sky130_fd_sc_hd__nor2_1 _10941_ (.A(_04844_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _10942_ (.A(net917),
    .B(net1983),
    .Y(_04847_));
 sky130_fd_sc_hd__and3_1 _10943_ (.A(net917),
    .B(net1983),
    .C(_04846_),
    .X(_04848_));
 sky130_fd_sc_hd__xnor2_1 _10944_ (.A(_04846_),
    .B(_04847_),
    .Y(_04849_));
 sky130_fd_sc_hd__a21o_1 _10945_ (.A1(_04811_),
    .A2(_04831_),
    .B1(_04842_),
    .X(_04850_));
 sky130_fd_sc_hd__nand3_1 _10946_ (.A(_04843_),
    .B(_04849_),
    .C(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(_04843_),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand3_1 _10948_ (.A(_04820_),
    .B(_04830_),
    .C(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__a21o_1 _10949_ (.A1(_04820_),
    .A2(_04830_),
    .B1(_04852_),
    .X(_04854_));
 sky130_fd_sc_hd__o211ai_2 _10950_ (.A1(_04845_),
    .A2(_04848_),
    .B1(_04853_),
    .C1(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__and2_1 _10951_ (.A(_04853_),
    .B(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__nor2_1 _10952_ (.A(_04829_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__xor2_1 _10953_ (.A(_04829_),
    .B(_04856_),
    .X(_04858_));
 sky130_fd_sc_hd__a211o_1 _10954_ (.A1(_04853_),
    .A2(_04854_),
    .B1(_04845_),
    .C1(_04848_),
    .X(_04859_));
 sky130_fd_sc_hd__a21o_1 _10955_ (.A1(_04843_),
    .A2(_04850_),
    .B1(_04849_),
    .X(_04860_));
 sky130_fd_sc_hd__a31o_1 _10956_ (.A1(_04835_),
    .A2(_04839_),
    .A3(_04840_),
    .B1(_04838_),
    .X(_04861_));
 sky130_fd_sc_hd__and4_1 _10957_ (.A(net69),
    .B(net917),
    .C(net1007),
    .D(net1010),
    .X(_04862_));
 sky130_fd_sc_hd__nand4_1 _10958_ (.A(net69),
    .B(net917),
    .C(net1007),
    .D(net1009),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2_1 _10959_ (.A(_04832_),
    .B(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _10960_ (.A(_04833_),
    .B(_04862_),
    .Y(_04865_));
 sky130_fd_sc_hd__a22oi_1 _10961_ (.A1(net1934),
    .A2(net992),
    .B1(net1970),
    .B2(net917),
    .Y(_04866_));
 sky130_fd_sc_hd__and4_1 _10962_ (.A(net917),
    .B(net1934),
    .C(net992),
    .D(net1970),
    .X(_04867_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(_04866_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _10964_ (.A(_04832_),
    .B(_04863_),
    .Y(_04869_));
 sky130_fd_sc_hd__a22o_1 _10965_ (.A1(net69),
    .A2(net1007),
    .B1(net1009),
    .B2(net953),
    .X(_04870_));
 sky130_fd_sc_hd__nand4_1 _10966_ (.A(_04865_),
    .B(_04868_),
    .C(_04869_),
    .D(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__a31o_1 _10967_ (.A1(_04868_),
    .A2(_04869_),
    .A3(_04870_),
    .B1(_04864_),
    .X(_04872_));
 sky130_fd_sc_hd__nand3_1 _10968_ (.A(_04841_),
    .B(_04861_),
    .C(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2_1 _10969_ (.A(net1615),
    .B(net1987),
    .Y(_04874_));
 sky130_fd_sc_hd__nand3_2 _10970_ (.A(net1615),
    .B(net1987),
    .C(_04867_),
    .Y(_04875_));
 sky130_fd_sc_hd__xnor2_1 _10971_ (.A(_04867_),
    .B(_04874_),
    .Y(_04876_));
 sky130_fd_sc_hd__and2_1 _10972_ (.A(net1934),
    .B(net1983),
    .X(_04877_));
 sky130_fd_sc_hd__or2_1 _10973_ (.A(_04876_),
    .B(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _10974_ (.A(_04876_),
    .B(_04877_),
    .Y(_04879_));
 sky130_fd_sc_hd__and2_1 _10975_ (.A(_04878_),
    .B(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__a21o_1 _10976_ (.A1(_04841_),
    .A2(_04861_),
    .B1(_04872_),
    .X(_04881_));
 sky130_fd_sc_hd__nand3_1 _10977_ (.A(_04873_),
    .B(_04880_),
    .C(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__a21bo_1 _10978_ (.A1(_04880_),
    .A2(_04881_),
    .B1_N(_04873_),
    .X(_04883_));
 sky130_fd_sc_hd__and3_2 _10979_ (.A(_04851_),
    .B(_04860_),
    .C(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__a21oi_2 _10980_ (.A1(_04851_),
    .A2(_04860_),
    .B1(_04883_),
    .Y(_04885_));
 sky130_fd_sc_hd__a211oi_4 _10981_ (.A1(_04875_),
    .A2(_04879_),
    .B1(_04884_),
    .C1(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__o211a_1 _10982_ (.A1(_04884_),
    .A2(_04886_),
    .B1(_04855_),
    .C1(_04859_),
    .X(_04887_));
 sky130_fd_sc_hd__a211o_1 _10983_ (.A1(_04855_),
    .A2(_04859_),
    .B1(_04884_),
    .C1(_04886_),
    .X(_04888_));
 sky130_fd_sc_hd__nand2b_1 _10984_ (.A_N(_04887_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__o211a_1 _10985_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04875_),
    .C1(_04879_),
    .X(_04890_));
 sky130_fd_sc_hd__a21o_1 _10986_ (.A1(_04873_),
    .A2(_04881_),
    .B1(_04880_),
    .X(_04891_));
 sky130_fd_sc_hd__a31o_1 _10987_ (.A1(_04865_),
    .A2(_04869_),
    .A3(_04870_),
    .B1(_04868_),
    .X(_04892_));
 sky130_fd_sc_hd__nand4_2 _10988_ (.A(net917),
    .B(net1934),
    .C(net1007),
    .D(net1010),
    .Y(_04893_));
 sky130_fd_sc_hd__nor2_1 _10989_ (.A(_04862_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__a22oi_1 _10990_ (.A1(net1615),
    .A2(net992),
    .B1(net1970),
    .B2(net1934),
    .Y(_04895_));
 sky130_fd_sc_hd__and4_1 _10991_ (.A(net1934),
    .B(net1615),
    .C(net992),
    .D(net1970),
    .X(_04896_));
 sky130_fd_sc_hd__nor2_1 _10992_ (.A(_04895_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_04862_),
    .B(_04893_),
    .Y(_04898_));
 sky130_fd_sc_hd__a22o_1 _10994_ (.A1(net917),
    .A2(net1007),
    .B1(net1010),
    .B2(net69),
    .X(_04899_));
 sky130_fd_sc_hd__and3b_1 _10995_ (.A_N(_04894_),
    .B(_04898_),
    .C(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__a31o_1 _10996_ (.A1(_04897_),
    .A2(_04898_),
    .A3(_04899_),
    .B1(_04894_),
    .X(_04901_));
 sky130_fd_sc_hd__and3_1 _10997_ (.A(_04871_),
    .B(_04892_),
    .C(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__a21o_1 _10998_ (.A1(net1615),
    .A2(net1983),
    .B1(_04896_),
    .X(_04903_));
 sky130_fd_sc_hd__nand2_1 _10999_ (.A(net1983),
    .B(_04896_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _11000_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21o_1 _11001_ (.A1(_04871_),
    .A2(_04892_),
    .B1(_04901_),
    .X(_04906_));
 sky130_fd_sc_hd__and2b_1 _11002_ (.A_N(_04902_),
    .B(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__a31o_1 _11003_ (.A1(_04903_),
    .A2(_04904_),
    .A3(_04906_),
    .B1(_04902_),
    .X(_04908_));
 sky130_fd_sc_hd__and3_1 _11004_ (.A(_04882_),
    .B(_04891_),
    .C(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__inv_2 _11005_ (.A(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__a21oi_1 _11006_ (.A1(_04882_),
    .A2(_04891_),
    .B1(_04908_),
    .Y(_04911_));
 sky130_fd_sc_hd__or3_2 _11007_ (.A(_04904_),
    .B(_04909_),
    .C(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__a211o_1 _11008_ (.A1(_04910_),
    .A2(_04912_),
    .B1(_04886_),
    .C1(_04890_),
    .X(_04913_));
 sky130_fd_sc_hd__xnor2_1 _11009_ (.A(_04905_),
    .B(_04907_),
    .Y(_04914_));
 sky130_fd_sc_hd__xnor2_1 _11010_ (.A(_04897_),
    .B(_04900_),
    .Y(_04915_));
 sky130_fd_sc_hd__and4_1 _11011_ (.A(net1934),
    .B(net1615),
    .C(net1007),
    .D(net1010),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _11012_ (.A(net1615),
    .B(net1970),
    .Y(_04917_));
 sky130_fd_sc_hd__a22oi_1 _11013_ (.A1(net1934),
    .A2(net1007),
    .B1(net1010),
    .B2(net917),
    .Y(_04918_));
 sky130_fd_sc_hd__a21oi_1 _11014_ (.A1(_04893_),
    .A2(_04916_),
    .B1(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__o21ai_1 _11015_ (.A1(_04893_),
    .A2(_04916_),
    .B1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__a2bb2o_1 _11016_ (.A1_N(_04917_),
    .A2_N(_04920_),
    .B1(_04893_),
    .B2(_04916_),
    .X(_04921_));
 sky130_fd_sc_hd__and2b_1 _11017_ (.A_N(_04915_),
    .B(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__and2_1 _11018_ (.A(_04914_),
    .B(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__o21ai_1 _11019_ (.A1(_04909_),
    .A2(_04911_),
    .B1(_04904_),
    .Y(_04924_));
 sky130_fd_sc_hd__and3_1 _11020_ (.A(_04912_),
    .B(_04923_),
    .C(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o211ai_2 _11021_ (.A1(_04886_),
    .A2(_04890_),
    .B1(_04910_),
    .C1(_04912_),
    .Y(_04926_));
 sky130_fd_sc_hd__and3_1 _11022_ (.A(_04913_),
    .B(_04925_),
    .C(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__a21bo_1 _11023_ (.A1(_04925_),
    .A2(_04926_),
    .B1_N(_04913_),
    .X(_04928_));
 sky130_fd_sc_hd__a21o_1 _11024_ (.A1(_04888_),
    .A2(_04928_),
    .B1(_04887_),
    .X(_04929_));
 sky130_fd_sc_hd__a21oi_1 _11025_ (.A1(_04858_),
    .A2(_04929_),
    .B1(_04857_),
    .Y(_04930_));
 sky130_fd_sc_hd__a211o_1 _11026_ (.A1(_04858_),
    .A2(_04929_),
    .B1(_04828_),
    .C1(_04857_),
    .X(_04931_));
 sky130_fd_sc_hd__and3_1 _11027_ (.A(_04798_),
    .B(_04827_),
    .C(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__a31o_1 _11028_ (.A1(_04798_),
    .A2(_04827_),
    .A3(_04931_),
    .B1(_04797_),
    .X(_04933_));
 sky130_fd_sc_hd__a311o_1 _11029_ (.A1(_04798_),
    .A2(_04827_),
    .A3(_04931_),
    .B1(_04797_),
    .C1(_04767_),
    .X(_04934_));
 sky130_fd_sc_hd__and3_1 _11030_ (.A(_04732_),
    .B(_04766_),
    .C(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a31o_1 _11031_ (.A1(_04732_),
    .A2(_04766_),
    .A3(_04934_),
    .B1(_04730_),
    .X(_04936_));
 sky130_fd_sc_hd__a21oi_2 _11032_ (.A1(_04701_),
    .A2(_04936_),
    .B1(_04699_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2b_1 _11033_ (.A_N(_04937_),
    .B(_04676_),
    .Y(_04938_));
 sky130_fd_sc_hd__xor2_2 _11034_ (.A(_04676_),
    .B(_04937_),
    .X(_04939_));
 sky130_fd_sc_hd__a22oi_1 _11035_ (.A1(net614),
    .A2(net2023),
    .B1(net717),
    .B2(net1407),
    .Y(_04940_));
 sky130_fd_sc_hd__and4_1 _11036_ (.A(net1407),
    .B(net614),
    .C(net2023),
    .D(net717),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _11037_ (.A(_04940_),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(net614),
    .B(net717),
    .Y(_04943_));
 sky130_fd_sc_hd__and4_1 _11039_ (.A(net614),
    .B(net2235),
    .C(net2023),
    .D(net2281),
    .X(_04944_));
 sky130_fd_sc_hd__a22o_1 _11040_ (.A1(net2235),
    .A2(net2023),
    .B1(net717),
    .B2(net614),
    .X(_04945_));
 sky130_fd_sc_hd__and2b_1 _11041_ (.A_N(_04944_),
    .B(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__nand2_1 _11042_ (.A(net1407),
    .B(net1821),
    .Y(_04947_));
 sky130_fd_sc_hd__a31o_1 _11043_ (.A1(net1407),
    .A2(net1821),
    .A3(_04945_),
    .B1(_04944_),
    .X(_04948_));
 sky130_fd_sc_hd__and2_1 _11044_ (.A(_04942_),
    .B(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__xor2_1 _11045_ (.A(_04946_),
    .B(_04947_),
    .X(_04950_));
 sky130_fd_sc_hd__nand4_1 _11046_ (.A(net2235),
    .B(net845),
    .C(net2023),
    .D(net717),
    .Y(_04951_));
 sky130_fd_sc_hd__a22o_1 _11047_ (.A1(net845),
    .A2(net2023),
    .B1(net717),
    .B2(net2235),
    .X(_04952_));
 sky130_fd_sc_hd__nand2_1 _11048_ (.A(_04951_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand2_1 _11049_ (.A(net614),
    .B(net1821),
    .Y(_04954_));
 sky130_fd_sc_hd__o21ai_1 _11050_ (.A1(_04953_),
    .A2(_04954_),
    .B1(_04951_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2b_2 _11051_ (.A_N(_04950_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__nor2_1 _11052_ (.A(_04942_),
    .B(_04948_),
    .Y(_04957_));
 sky130_fd_sc_hd__or2_2 _11053_ (.A(_04949_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__o21bai_4 _11054_ (.A1(_04956_),
    .A2(_04958_),
    .B1_N(_04949_),
    .Y(_04959_));
 sky130_fd_sc_hd__and3_2 _11055_ (.A(net1407),
    .B(net2023),
    .C(_04943_),
    .X(_04960_));
 sky130_fd_sc_hd__xnor2_4 _11056_ (.A(_04959_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__inv_2 _11057_ (.A(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__nand2b_1 _11058_ (.A_N(_04955_),
    .B(_04950_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_04956_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__xnor2_1 _11060_ (.A(_04953_),
    .B(_04954_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand4_1 _11061_ (.A(net845),
    .B(net1001),
    .C(net2023),
    .D(net717),
    .Y(_04966_));
 sky130_fd_sc_hd__a22o_1 _11062_ (.A1(net1001),
    .A2(net2023),
    .B1(net717),
    .B2(net845),
    .X(_04967_));
 sky130_fd_sc_hd__nand2_1 _11063_ (.A(_04966_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__nand2_1 _11064_ (.A(net2235),
    .B(net1821),
    .Y(_04969_));
 sky130_fd_sc_hd__o21ai_1 _11065_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_04966_),
    .Y(_04970_));
 sky130_fd_sc_hd__and2b_1 _11066_ (.A_N(_04965_),
    .B(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__and2b_1 _11067_ (.A_N(_04970_),
    .B(_04965_),
    .X(_04972_));
 sky130_fd_sc_hd__nor2_1 _11068_ (.A(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_1 _11069_ (.A(net1407),
    .B(net782),
    .Y(_04974_));
 sky130_fd_sc_hd__a31oi_1 _11070_ (.A1(net1407),
    .A2(net782),
    .A3(_04973_),
    .B1(_04971_),
    .Y(_04975_));
 sky130_fd_sc_hd__or2_1 _11071_ (.A(_04964_),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__nor2_2 _11072_ (.A(_04958_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__xnor2_4 _11073_ (.A(_04961_),
    .B(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand2_1 _11074_ (.A(_04964_),
    .B(_04975_),
    .Y(_04979_));
 sky130_fd_sc_hd__and2_1 _11075_ (.A(_04976_),
    .B(_04979_),
    .X(_04980_));
 sky130_fd_sc_hd__xnor2_1 _11076_ (.A(_04973_),
    .B(_04974_),
    .Y(_04981_));
 sky130_fd_sc_hd__xnor2_1 _11077_ (.A(_04968_),
    .B(_04969_),
    .Y(_04982_));
 sky130_fd_sc_hd__and4_1 _11078_ (.A(net1001),
    .B(net965),
    .C(net2023),
    .D(net717),
    .X(_04983_));
 sky130_fd_sc_hd__a22o_1 _11079_ (.A1(net965),
    .A2(net2023),
    .B1(net717),
    .B2(net1001),
    .X(_04984_));
 sky130_fd_sc_hd__nand2b_1 _11080_ (.A_N(_04983_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _11081_ (.A(net845),
    .B(net1821),
    .Y(_04986_));
 sky130_fd_sc_hd__a31o_1 _11082_ (.A1(net845),
    .A2(net1821),
    .A3(_04984_),
    .B1(_04983_),
    .X(_04987_));
 sky130_fd_sc_hd__and2b_1 _11083_ (.A_N(_04982_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__xor2_1 _11084_ (.A(_04982_),
    .B(_04987_),
    .X(_04989_));
 sky130_fd_sc_hd__a22oi_1 _11085_ (.A1(net614),
    .A2(net782),
    .B1(net1004),
    .B2(net1407),
    .Y(_04990_));
 sky130_fd_sc_hd__and4_1 _11086_ (.A(net1407),
    .B(net614),
    .C(net782),
    .D(net1004),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _11087_ (.A(_04990_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__and2b_1 _11088_ (.A_N(_04989_),
    .B(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__o21a_1 _11089_ (.A1(_04988_),
    .A2(_04993_),
    .B1(_04981_),
    .X(_04994_));
 sky130_fd_sc_hd__or3_1 _11090_ (.A(_04981_),
    .B(_04988_),
    .C(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__and2b_1 _11091_ (.A_N(_04994_),
    .B(_04995_),
    .X(_04996_));
 sky130_fd_sc_hd__a21oi_1 _11092_ (.A1(_04991_),
    .A2(_04995_),
    .B1(_04994_),
    .Y(_04997_));
 sky130_fd_sc_hd__and2b_1 _11093_ (.A_N(_04997_),
    .B(_04980_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(_04956_),
    .B(_04976_),
    .Y(_04999_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(_04958_),
    .B(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _11096_ (.A(_04998_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__or2_1 _11097_ (.A(_04998_),
    .B(_05000_),
    .X(_05002_));
 sky130_fd_sc_hd__nand2_2 _11098_ (.A(_05001_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__and2b_1 _11099_ (.A_N(_04980_),
    .B(_04997_),
    .X(_05004_));
 sky130_fd_sc_hd__or2_1 _11100_ (.A(_04998_),
    .B(_05004_),
    .X(_05005_));
 sky130_fd_sc_hd__xnor2_1 _11101_ (.A(_04991_),
    .B(_04996_),
    .Y(_05006_));
 sky130_fd_sc_hd__xnor2_1 _11102_ (.A(_04989_),
    .B(_04992_),
    .Y(_05007_));
 sky130_fd_sc_hd__xnor2_1 _11103_ (.A(_04985_),
    .B(_04986_),
    .Y(_05008_));
 sky130_fd_sc_hd__nand4_2 _11104_ (.A(net965),
    .B(net968),
    .C(net2023),
    .D(net2281),
    .Y(_05009_));
 sky130_fd_sc_hd__a22o_1 _11105_ (.A1(net968),
    .A2(net2023),
    .B1(net717),
    .B2(net965),
    .X(_05010_));
 sky130_fd_sc_hd__nand4_1 _11106_ (.A(net1001),
    .B(net1821),
    .C(_05009_),
    .D(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _11107_ (.A(_05009_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__and2b_1 _11108_ (.A_N(_05008_),
    .B(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a22o_1 _11109_ (.A1(net2235),
    .A2(net782),
    .B1(net1004),
    .B2(net614),
    .X(_05014_));
 sky130_fd_sc_hd__and4_1 _11110_ (.A(net614),
    .B(net2235),
    .C(net782),
    .D(net1004),
    .X(_05015_));
 sky130_fd_sc_hd__nand4_1 _11111_ (.A(net614),
    .B(net2235),
    .C(net781),
    .D(net1004),
    .Y(_05016_));
 sky130_fd_sc_hd__a22oi_1 _11112_ (.A1(net1407),
    .A2(net788),
    .B1(_05014_),
    .B2(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__and4_1 _11113_ (.A(net1407),
    .B(net788),
    .C(_05014_),
    .D(_05016_),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _11114_ (.A(_05017_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__xor2_1 _11115_ (.A(_05008_),
    .B(_05012_),
    .X(_05020_));
 sky130_fd_sc_hd__nor2_1 _11116_ (.A(_05019_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__o21ai_2 _11117_ (.A1(_05013_),
    .A2(_05021_),
    .B1(_05007_),
    .Y(_05022_));
 sky130_fd_sc_hd__or3_2 _11118_ (.A(_05007_),
    .B(_05013_),
    .C(_05021_),
    .X(_05023_));
 sky130_fd_sc_hd__o211ai_4 _11119_ (.A1(_05015_),
    .A2(_05018_),
    .B1(_05022_),
    .C1(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _11120_ (.A(_05022_),
    .B(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2b_1 _11121_ (.A_N(_05006_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nor2_1 _11122_ (.A(_05005_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__and2_1 _11123_ (.A(_05005_),
    .B(_05026_),
    .X(_05028_));
 sky130_fd_sc_hd__nor2_1 _11124_ (.A(_05027_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__xor2_1 _11125_ (.A(_05006_),
    .B(_05025_),
    .X(_05030_));
 sky130_fd_sc_hd__a211o_1 _11126_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_05015_),
    .C1(_05018_),
    .X(_05031_));
 sky130_fd_sc_hd__xor2_1 _11127_ (.A(_05019_),
    .B(_05020_),
    .X(_05032_));
 sky130_fd_sc_hd__a22o_1 _11128_ (.A1(net1001),
    .A2(net1821),
    .B1(_05009_),
    .B2(_05010_),
    .X(_05033_));
 sky130_fd_sc_hd__nand4_2 _11129_ (.A(net968),
    .B(net1626),
    .C(net2023),
    .D(net717),
    .Y(_05034_));
 sky130_fd_sc_hd__and2_1 _11130_ (.A(net965),
    .B(net1821),
    .X(_05035_));
 sky130_fd_sc_hd__a22o_1 _11131_ (.A1(net1626),
    .A2(net2023),
    .B1(net717),
    .B2(net968),
    .X(_05036_));
 sky130_fd_sc_hd__nand3_1 _11132_ (.A(_05034_),
    .B(_05035_),
    .C(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21bo_1 _11133_ (.A1(_05035_),
    .A2(_05036_),
    .B1_N(_05034_),
    .X(_05038_));
 sky130_fd_sc_hd__and3_1 _11134_ (.A(_05011_),
    .B(_05033_),
    .C(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__a22oi_2 _11135_ (.A1(net845),
    .A2(net781),
    .B1(net1003),
    .B2(net2235),
    .Y(_05040_));
 sky130_fd_sc_hd__and4_1 _11136_ (.A(net2235),
    .B(net845),
    .C(net781),
    .D(net1003),
    .X(_05041_));
 sky130_fd_sc_hd__nor2_1 _11137_ (.A(_05040_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _11138_ (.A(net1508),
    .B(net788),
    .Y(_05043_));
 sky130_fd_sc_hd__xnor2_1 _11139_ (.A(_05042_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__a21oi_1 _11140_ (.A1(_05011_),
    .A2(_05033_),
    .B1(_05038_),
    .Y(_05045_));
 sky130_fd_sc_hd__or3b_1 _11141_ (.A(_05039_),
    .B(_05045_),
    .C_N(_05044_),
    .X(_05046_));
 sky130_fd_sc_hd__and2b_1 _11142_ (.A_N(_05039_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__and2b_1 _11143_ (.A_N(_05047_),
    .B(_05032_),
    .X(_05048_));
 sky130_fd_sc_hd__o21ba_1 _11144_ (.A1(_05040_),
    .A2(_05043_),
    .B1_N(_05041_),
    .X(_05049_));
 sky130_fd_sc_hd__xnor2_1 _11145_ (.A(_05032_),
    .B(_05047_),
    .Y(_05050_));
 sky130_fd_sc_hd__and2b_1 _11146_ (.A_N(_05049_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__o211ai_4 _11147_ (.A1(_05048_),
    .A2(_05051_),
    .B1(_05024_),
    .C1(_05031_),
    .Y(_05052_));
 sky130_fd_sc_hd__a211o_1 _11148_ (.A1(_05024_),
    .A2(_05031_),
    .B1(_05048_),
    .C1(_05051_),
    .X(_05053_));
 sky130_fd_sc_hd__nand2_1 _11149_ (.A(_05052_),
    .B(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__xnor2_1 _11150_ (.A(_05049_),
    .B(_05050_),
    .Y(_05055_));
 sky130_fd_sc_hd__o21bai_1 _11151_ (.A1(_05039_),
    .A2(_05045_),
    .B1_N(_05044_),
    .Y(_05056_));
 sky130_fd_sc_hd__a21o_1 _11152_ (.A1(_05034_),
    .A2(_05036_),
    .B1(_05035_),
    .X(_05057_));
 sky130_fd_sc_hd__and4_1 _11153_ (.A(net968),
    .B(net1626),
    .C(net717),
    .D(net1821),
    .X(_05058_));
 sky130_fd_sc_hd__inv_2 _11154_ (.A(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand3_1 _11155_ (.A(_05037_),
    .B(_05057_),
    .C(_05058_),
    .Y(_05060_));
 sky130_fd_sc_hd__a22oi_2 _11156_ (.A1(net1001),
    .A2(net781),
    .B1(net3710),
    .B2(net2437),
    .Y(_05061_));
 sky130_fd_sc_hd__and4_1 _11157_ (.A(net2437),
    .B(net2442),
    .C(net781),
    .D(net3710),
    .X(_05062_));
 sky130_fd_sc_hd__nor2_1 _11158_ (.A(_05061_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _11159_ (.A(net2235),
    .B(net788),
    .Y(_05064_));
 sky130_fd_sc_hd__xnor2_1 _11160_ (.A(_05063_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__a21o_1 _11161_ (.A1(_05037_),
    .A2(_05057_),
    .B1(_05058_),
    .X(_05066_));
 sky130_fd_sc_hd__nand3_1 _11162_ (.A(_05060_),
    .B(_05065_),
    .C(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__a21bo_1 _11163_ (.A1(_05065_),
    .A2(_05066_),
    .B1_N(_05060_),
    .X(_05068_));
 sky130_fd_sc_hd__and3_1 _11164_ (.A(_05046_),
    .B(_05056_),
    .C(_05068_),
    .X(_05069_));
 sky130_fd_sc_hd__o21ba_1 _11165_ (.A1(net3711),
    .A2(_05064_),
    .B1_N(_05062_),
    .X(_05070_));
 sky130_fd_sc_hd__nand2_1 _11166_ (.A(net1407),
    .B(net1954),
    .Y(_05071_));
 sky130_fd_sc_hd__nor2_1 _11167_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__xnor2_1 _11168_ (.A(_05070_),
    .B(_05071_),
    .Y(_05073_));
 sky130_fd_sc_hd__a21oi_1 _11169_ (.A1(_05046_),
    .A2(_05056_),
    .B1(_05068_),
    .Y(_05074_));
 sky130_fd_sc_hd__nor3_1 _11170_ (.A(_05069_),
    .B(_05073_),
    .C(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _11171_ (.A(_05069_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__and2b_1 _11172_ (.A_N(_05076_),
    .B(_05055_),
    .X(_05077_));
 sky130_fd_sc_hd__xnor2_1 _11173_ (.A(_05055_),
    .B(_05076_),
    .Y(_05078_));
 sky130_fd_sc_hd__and2_1 _11174_ (.A(_05072_),
    .B(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__or2_1 _11175_ (.A(_05077_),
    .B(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__and3_1 _11176_ (.A(_05052_),
    .B(_05053_),
    .C(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__o21bai_1 _11177_ (.A1(_05077_),
    .A2(_05079_),
    .B1_N(_05054_),
    .Y(_05082_));
 sky130_fd_sc_hd__a21oi_1 _11178_ (.A1(_05052_),
    .A2(_05082_),
    .B1(_05030_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _11179_ (.A(_05030_),
    .B(_05052_),
    .Y(_05084_));
 sky130_fd_sc_hd__xnor2_2 _11180_ (.A(_05054_),
    .B(_05080_),
    .Y(_05085_));
 sky130_fd_sc_hd__xnor2_1 _11181_ (.A(_05072_),
    .B(_05078_),
    .Y(_05086_));
 sky130_fd_sc_hd__o21a_1 _11182_ (.A1(_05069_),
    .A2(_05074_),
    .B1(_05073_),
    .X(_05087_));
 sky130_fd_sc_hd__or2_2 _11183_ (.A(_05075_),
    .B(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__a21o_1 _11184_ (.A1(_05060_),
    .A2(_05066_),
    .B1(_05065_),
    .X(_05089_));
 sky130_fd_sc_hd__and4_1 _11185_ (.A(net2442),
    .B(net3600),
    .C(net782),
    .D(net1004),
    .X(_05090_));
 sky130_fd_sc_hd__nand4_2 _11186_ (.A(net2442),
    .B(net965),
    .C(net782),
    .D(net1004),
    .Y(_05091_));
 sky130_fd_sc_hd__a22o_1 _11187_ (.A1(net3600),
    .A2(net782),
    .B1(net1004),
    .B2(net1001),
    .X(_05092_));
 sky130_fd_sc_hd__and4_1 _11188_ (.A(net845),
    .B(net2297),
    .C(_05091_),
    .D(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__nand4_1 _11189_ (.A(net845),
    .B(net788),
    .C(_05091_),
    .D(_05092_),
    .Y(_05094_));
 sky130_fd_sc_hd__a22o_1 _11190_ (.A1(net845),
    .A2(net788),
    .B1(_05091_),
    .B2(_05092_),
    .X(_05095_));
 sky130_fd_sc_hd__a22o_1 _11191_ (.A1(net1626),
    .A2(net717),
    .B1(net1821),
    .B2(net968),
    .X(_05096_));
 sky130_fd_sc_hd__nand4_2 _11192_ (.A(_05059_),
    .B(_05094_),
    .C(_05095_),
    .D(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand3b_2 _11193_ (.A_N(_05097_),
    .B(_05089_),
    .C(_05067_),
    .Y(_05098_));
 sky130_fd_sc_hd__o211a_1 _11194_ (.A1(_05090_),
    .A2(_05093_),
    .B1(net614),
    .C1(net1954),
    .X(_05099_));
 sky130_fd_sc_hd__a211oi_1 _11195_ (.A1(net614),
    .A2(net1954),
    .B1(_05090_),
    .C1(_05093_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_1 _11196_ (.A(_05099_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(net1407),
    .B(net2333),
    .Y(_05102_));
 sky130_fd_sc_hd__xnor2_1 _11198_ (.A(_05101_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__a21bo_1 _11199_ (.A1(_05067_),
    .A2(_05089_),
    .B1_N(_05097_),
    .X(_05104_));
 sky130_fd_sc_hd__nand3_2 _11200_ (.A(_05098_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2_2 _11201_ (.A(_05098_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2b_1 _11202_ (.A_N(_05088_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__a31o_2 _11203_ (.A1(net1407),
    .A2(net2333),
    .A3(_05101_),
    .B1(_05099_),
    .X(_05108_));
 sky130_fd_sc_hd__xnor2_4 _11204_ (.A(_05088_),
    .B(_05106_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand2_1 _11205_ (.A(_05108_),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__and3_1 _11206_ (.A(_05086_),
    .B(_05107_),
    .C(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__nand3_2 _11207_ (.A(_05086_),
    .B(_05107_),
    .C(_05110_),
    .Y(_05112_));
 sky130_fd_sc_hd__a21oi_1 _11208_ (.A1(_05107_),
    .A2(_05110_),
    .B1(_05086_),
    .Y(_05113_));
 sky130_fd_sc_hd__xnor2_4 _11209_ (.A(_05108_),
    .B(_05109_),
    .Y(_05114_));
 sky130_fd_sc_hd__a21o_1 _11210_ (.A1(_05098_),
    .A2(_05104_),
    .B1(_05103_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _11211_ (.A1(_05094_),
    .A2(_05095_),
    .B1(_05096_),
    .B2(_05059_),
    .X(_05116_));
 sky130_fd_sc_hd__nand2_1 _11212_ (.A(net1626),
    .B(net1821),
    .Y(_05117_));
 sky130_fd_sc_hd__and4_1 _11213_ (.A(net965),
    .B(net968),
    .C(net782),
    .D(net1004),
    .X(_05118_));
 sky130_fd_sc_hd__a22oi_1 _11214_ (.A1(net3676),
    .A2(net782),
    .B1(net1004),
    .B2(net965),
    .Y(_05119_));
 sky130_fd_sc_hd__a22o_1 _11215_ (.A1(net3676),
    .A2(net782),
    .B1(net1004),
    .B2(net965),
    .X(_05120_));
 sky130_fd_sc_hd__and4b_1 _11216_ (.A_N(_05118_),
    .B(_05120_),
    .C(net1001),
    .D(net788),
    .X(_05121_));
 sky130_fd_sc_hd__o2bb2a_1 _11217_ (.A1_N(net1001),
    .A2_N(net788),
    .B1(_05118_),
    .B2(_05119_),
    .X(_05122_));
 sky130_fd_sc_hd__nor3_1 _11218_ (.A(_05117_),
    .B(_05121_),
    .C(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__and3_1 _11219_ (.A(_05097_),
    .B(_05116_),
    .C(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__nand3_1 _11220_ (.A(_05097_),
    .B(_05116_),
    .C(_05123_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_1 _11221_ (.A(net614),
    .B(net809),
    .Y(_05126_));
 sky130_fd_sc_hd__a31o_1 _11222_ (.A1(net1001),
    .A2(net788),
    .A3(_05120_),
    .B1(_05118_),
    .X(_05127_));
 sky130_fd_sc_hd__nand2_1 _11223_ (.A(net2235),
    .B(net1954),
    .Y(_05128_));
 sky130_fd_sc_hd__and3_1 _11224_ (.A(net2235),
    .B(net1954),
    .C(_05127_),
    .X(_05129_));
 sky130_fd_sc_hd__xnor2_1 _11225_ (.A(_05127_),
    .B(_05128_),
    .Y(_05130_));
 sky130_fd_sc_hd__and3_1 _11226_ (.A(net614),
    .B(net2333),
    .C(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__xnor2_1 _11227_ (.A(_05126_),
    .B(_05130_),
    .Y(_05132_));
 sky130_fd_sc_hd__a21o_1 _11228_ (.A1(_05097_),
    .A2(_05116_),
    .B1(_05123_),
    .X(_05133_));
 sky130_fd_sc_hd__and3_2 _11229_ (.A(_05125_),
    .B(_05132_),
    .C(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__o211ai_4 _11230_ (.A1(_05124_),
    .A2(_05134_),
    .B1(_05105_),
    .C1(_05115_),
    .Y(_05135_));
 sky130_fd_sc_hd__a211o_1 _11231_ (.A1(_05105_),
    .A2(_05115_),
    .B1(_05124_),
    .C1(_05134_),
    .X(_05136_));
 sky130_fd_sc_hd__o211ai_2 _11232_ (.A1(net3173),
    .A2(_05131_),
    .B1(_05135_),
    .C1(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_2 _11233_ (.A(_05135_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__and2b_1 _11234_ (.A_N(_05114_),
    .B(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__a211o_1 _11235_ (.A1(_05135_),
    .A2(_05136_),
    .B1(net3173),
    .C1(_05131_),
    .X(_05140_));
 sky130_fd_sc_hd__a21oi_1 _11236_ (.A1(_05125_),
    .A2(_05133_),
    .B1(_05132_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(net2235),
    .B(net2333),
    .Y(_05142_));
 sky130_fd_sc_hd__and3_1 _11238_ (.A(net968),
    .B(net1626),
    .C(net1004),
    .X(_05143_));
 sky130_fd_sc_hd__nand2_1 _11239_ (.A(net965),
    .B(net788),
    .Y(_05144_));
 sky130_fd_sc_hd__a22o_1 _11240_ (.A1(net1626),
    .A2(net782),
    .B1(net1004),
    .B2(net968),
    .X(_05145_));
 sky130_fd_sc_hd__a21bo_1 _11241_ (.A1(net782),
    .A2(_05143_),
    .B1_N(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__a32o_1 _11242_ (.A1(net965),
    .A2(net788),
    .A3(_05145_),
    .B1(_05143_),
    .B2(net782),
    .X(_05147_));
 sky130_fd_sc_hd__nand2_1 _11243_ (.A(net845),
    .B(net1954),
    .Y(_05148_));
 sky130_fd_sc_hd__and3_1 _11244_ (.A(net845),
    .B(net1954),
    .C(_05147_),
    .X(_05149_));
 sky130_fd_sc_hd__xnor2_1 _11245_ (.A(_05147_),
    .B(_05148_),
    .Y(_05150_));
 sky130_fd_sc_hd__xnor2_1 _11246_ (.A(_05142_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21a_1 _11247_ (.A1(_05121_),
    .A2(_05122_),
    .B1(_05117_),
    .X(_05152_));
 sky130_fd_sc_hd__nor2_1 _11248_ (.A(_05123_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(_05151_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__nor3_2 _11250_ (.A(_05134_),
    .B(_05141_),
    .C(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__a31o_1 _11251_ (.A1(net2235),
    .A2(net2333),
    .A3(_05150_),
    .B1(_05149_),
    .X(_05156_));
 sky130_fd_sc_hd__inv_2 _11252_ (.A(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__o21a_1 _11253_ (.A1(_05134_),
    .A2(_05141_),
    .B1(_05154_),
    .X(_05158_));
 sky130_fd_sc_hd__nor3_1 _11254_ (.A(_05155_),
    .B(_05157_),
    .C(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__or3_1 _11255_ (.A(_05155_),
    .B(_05157_),
    .C(_05158_),
    .X(_05160_));
 sky130_fd_sc_hd__o211a_1 _11256_ (.A1(_05155_),
    .A2(_05159_),
    .B1(_05137_),
    .C1(_05140_),
    .X(_05161_));
 sky130_fd_sc_hd__a211o_1 _11257_ (.A1(_05137_),
    .A2(_05140_),
    .B1(_05155_),
    .C1(_05159_),
    .X(_05162_));
 sky130_fd_sc_hd__o21ai_1 _11258_ (.A1(_05155_),
    .A2(_05158_),
    .B1(_05157_),
    .Y(_05163_));
 sky130_fd_sc_hd__xnor2_1 _11259_ (.A(_05151_),
    .B(_05153_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _11260_ (.A(net845),
    .B(net809),
    .Y(_05165_));
 sky130_fd_sc_hd__and4_1 _11261_ (.A(net968),
    .B(net1626),
    .C(net1004),
    .D(net788),
    .X(_05166_));
 sky130_fd_sc_hd__inv_2 _11262_ (.A(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__a21oi_1 _11263_ (.A1(net1001),
    .A2(net1954),
    .B1(_05166_),
    .Y(_05168_));
 sky130_fd_sc_hd__and3_1 _11264_ (.A(net1001),
    .B(net1954),
    .C(_05166_),
    .X(_05169_));
 sky130_fd_sc_hd__nor2_1 _11265_ (.A(_05168_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__xnor2_1 _11266_ (.A(_05165_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__xor2_1 _11267_ (.A(_05144_),
    .B(_05146_),
    .X(_05172_));
 sky130_fd_sc_hd__nand2_1 _11268_ (.A(_05171_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__nor2_1 _11269_ (.A(_05164_),
    .B(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__a31o_1 _11270_ (.A1(net845),
    .A2(net3623),
    .A3(_05170_),
    .B1(_05169_),
    .X(_05175_));
 sky130_fd_sc_hd__xor2_1 _11271_ (.A(_05164_),
    .B(_05173_),
    .X(_05176_));
 sky130_fd_sc_hd__and2_1 _11272_ (.A(_05175_),
    .B(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__o211a_1 _11273_ (.A1(_05174_),
    .A2(_05177_),
    .B1(_05160_),
    .C1(_05163_),
    .X(_05178_));
 sky130_fd_sc_hd__a211o_1 _11274_ (.A1(_05160_),
    .A2(_05163_),
    .B1(_05174_),
    .C1(_05177_),
    .X(_05179_));
 sky130_fd_sc_hd__and2b_1 _11275_ (.A_N(_05178_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__xnor2_1 _11276_ (.A(_05175_),
    .B(_05176_),
    .Y(_05181_));
 sky130_fd_sc_hd__xnor2_1 _11277_ (.A(_05171_),
    .B(_05172_),
    .Y(_05182_));
 sky130_fd_sc_hd__and4_1 _11278_ (.A(net1001),
    .B(net965),
    .C(net1954),
    .D(net809),
    .X(_05183_));
 sky130_fd_sc_hd__inv_2 _11279_ (.A(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__a22o_1 _11280_ (.A1(net1626),
    .A2(net1004),
    .B1(net788),
    .B2(net968),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_1 _11281_ (.A1(net965),
    .A2(net1954),
    .B1(net809),
    .B2(net1001),
    .X(_05186_));
 sky130_fd_sc_hd__or4bb_1 _11282_ (.A(_05166_),
    .B(_05183_),
    .C_N(_05185_),
    .D_N(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _11283_ (.A(_05184_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand2b_1 _11284_ (.A_N(_05182_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__xor2_1 _11285_ (.A(_05182_),
    .B(_05188_),
    .X(_05190_));
 sky130_fd_sc_hd__a22o_1 _11286_ (.A1(_05167_),
    .A2(_05185_),
    .B1(_05186_),
    .B2(_05184_),
    .X(_05191_));
 sky130_fd_sc_hd__and4_1 _11287_ (.A(net965),
    .B(net968),
    .C(net1954),
    .D(net809),
    .X(_05192_));
 sky130_fd_sc_hd__a22o_1 _11288_ (.A1(net968),
    .A2(net1954),
    .B1(net2333),
    .B2(net965),
    .X(_05193_));
 sky130_fd_sc_hd__inv_2 _11289_ (.A(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__and4b_1 _11290_ (.A_N(_05192_),
    .B(_05193_),
    .C(net1626),
    .D(net2298),
    .X(_05195_));
 sky130_fd_sc_hd__or2_1 _11291_ (.A(_05192_),
    .B(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__and3_1 _11292_ (.A(_05187_),
    .B(_05191_),
    .C(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__o2bb2a_1 _11293_ (.A1_N(net1626),
    .A2_N(net2298),
    .B1(_05192_),
    .B2(_05194_),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_1 _11294_ (.A(_05195_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__and4_1 _11295_ (.A(net968),
    .B(net1626),
    .C(net1954),
    .D(net2333),
    .X(_05200_));
 sky130_fd_sc_hd__inv_2 _11296_ (.A(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__and2_1 _11297_ (.A(_05199_),
    .B(_05200_),
    .X(_05202_));
 sky130_fd_sc_hd__a21oi_1 _11298_ (.A1(_05187_),
    .A2(_05191_),
    .B1(_05196_),
    .Y(_05203_));
 sky130_fd_sc_hd__nor2_1 _11299_ (.A(_05197_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__a21oi_1 _11300_ (.A1(_05202_),
    .A2(_05204_),
    .B1(_05197_),
    .Y(_05205_));
 sky130_fd_sc_hd__or2_1 _11301_ (.A(_05190_),
    .B(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__a21oi_2 _11302_ (.A1(_05189_),
    .A2(_05206_),
    .B1(_05181_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21o_1 _11303_ (.A1(_05179_),
    .A2(_05207_),
    .B1(_05178_),
    .X(_05208_));
 sky130_fd_sc_hd__a21o_2 _11304_ (.A1(_05162_),
    .A2(_05208_),
    .B1(_05161_),
    .X(_05209_));
 sky130_fd_sc_hd__xnor2_4 _11305_ (.A(_05114_),
    .B(_05138_),
    .Y(_05210_));
 sky130_fd_sc_hd__a21o_1 _11306_ (.A1(_05209_),
    .A2(_05210_),
    .B1(_05139_),
    .X(_05211_));
 sky130_fd_sc_hd__a211o_1 _11307_ (.A1(_05209_),
    .A2(_05210_),
    .B1(_05113_),
    .C1(_05139_),
    .X(_05212_));
 sky130_fd_sc_hd__and3_1 _11308_ (.A(_05085_),
    .B(_05112_),
    .C(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__a41o_1 _11309_ (.A1(_05084_),
    .A2(_05085_),
    .A3(_05112_),
    .A4(_05212_),
    .B1(_05083_),
    .X(_05214_));
 sky130_fd_sc_hd__a21oi_2 _11310_ (.A1(_05029_),
    .A2(_05214_),
    .B1(_05027_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21a_2 _11311_ (.A1(_05003_),
    .A2(_05215_),
    .B1(_05001_),
    .X(_05216_));
 sky130_fd_sc_hd__and2b_1 _11312_ (.A_N(_05216_),
    .B(_04978_),
    .X(_05217_));
 sky130_fd_sc_hd__xor2_4 _11313_ (.A(_04978_),
    .B(_05216_),
    .X(_05218_));
 sky130_fd_sc_hd__or2_1 _11314_ (.A(_04939_),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__xnor2_2 _11315_ (.A(_04939_),
    .B(_05218_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand4_4 _11316_ (.A(net1421),
    .B(net1156),
    .C(net1837),
    .D(net872),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _11317_ (.A(net1471),
    .B(net1837),
    .Y(_05222_));
 sky130_fd_sc_hd__nand2_1 _11318_ (.A(net1421),
    .B(net714),
    .Y(_05223_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(net714),
    .A1(_05223_),
    .S(_05221_),
    .X(_05224_));
 sky130_fd_sc_hd__o22a_1 _11320_ (.A1(_00665_),
    .A2(_05221_),
    .B1(_05222_),
    .B2(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__and3_1 _11321_ (.A(net1421),
    .B(net1837),
    .C(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__xor2_1 _11322_ (.A(_05222_),
    .B(_05224_),
    .X(_05227_));
 sky130_fd_sc_hd__and4_1 _11323_ (.A(net1421),
    .B(net1995),
    .C(net1837),
    .D(net2003),
    .X(_05228_));
 sky130_fd_sc_hd__a22oi_1 _11324_ (.A1(net1995),
    .A2(net1837),
    .B1(net2003),
    .B2(net1421),
    .Y(_05229_));
 sky130_fd_sc_hd__and4bb_1 _11325_ (.A_N(_05228_),
    .B_N(_05229_),
    .C(net1471),
    .D(net872),
    .X(_05230_));
 sky130_fd_sc_hd__or2_1 _11326_ (.A(_05228_),
    .B(_05230_),
    .X(_05231_));
 sky130_fd_sc_hd__and3_1 _11327_ (.A(net1471),
    .B(net714),
    .C(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__a22o_1 _11328_ (.A1(net1156),
    .A2(net1837),
    .B1(net872),
    .B2(net1421),
    .X(_05233_));
 sky130_fd_sc_hd__a21oi_1 _11329_ (.A1(net1471),
    .A2(net714),
    .B1(_05231_),
    .Y(_05234_));
 sky130_fd_sc_hd__nor2_1 _11330_ (.A(_05232_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__and3_1 _11331_ (.A(_05221_),
    .B(_05233_),
    .C(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__o21a_1 _11332_ (.A1(_05232_),
    .A2(_05236_),
    .B1(_05227_),
    .X(_05237_));
 sky130_fd_sc_hd__and2_1 _11333_ (.A(_05226_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__nor2_1 _11334_ (.A(_05226_),
    .B(_05237_),
    .Y(_05239_));
 sky130_fd_sc_hd__or2_2 _11335_ (.A(_05238_),
    .B(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__a21oi_1 _11336_ (.A1(_05221_),
    .A2(_05233_),
    .B1(_05235_),
    .Y(_05241_));
 sky130_fd_sc_hd__or2_1 _11337_ (.A(_05236_),
    .B(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__o2bb2a_1 _11338_ (.A1_N(net1471),
    .A2_N(net872),
    .B1(_05228_),
    .B2(_05229_),
    .X(_05243_));
 sky130_fd_sc_hd__or2_1 _11339_ (.A(_05230_),
    .B(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__a22oi_1 _11340_ (.A1(net2243),
    .A2(net1837),
    .B1(net2003),
    .B2(net1471),
    .Y(_05245_));
 sky130_fd_sc_hd__and4_1 _11341_ (.A(net1471),
    .B(net2243),
    .C(net1837),
    .D(net2003),
    .X(_05246_));
 sky130_fd_sc_hd__nor2_1 _11342_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__a21oi_1 _11343_ (.A1(net1156),
    .A2(net872),
    .B1(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__and3_1 _11344_ (.A(net1156),
    .B(net872),
    .C(_05247_),
    .X(_05249_));
 sky130_fd_sc_hd__nor2_1 _11345_ (.A(_05248_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_1 _11346_ (.A(net1471),
    .B(net935),
    .Y(_05251_));
 sky130_fd_sc_hd__and3_1 _11347_ (.A(net1421),
    .B(net1668),
    .C(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__and4_1 _11348_ (.A(net1421),
    .B(net1471),
    .C(net1668),
    .D(net935),
    .X(_05253_));
 sky130_fd_sc_hd__a21oi_2 _11349_ (.A1(_05250_),
    .A2(_05252_),
    .B1(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__xnor2_2 _11350_ (.A(_05244_),
    .B(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__nor2_1 _11351_ (.A(_05246_),
    .B(_05249_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_1 _11352_ (.A(net1156),
    .B(net714),
    .Y(_05257_));
 sky130_fd_sc_hd__or2_1 _11353_ (.A(_05256_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xnor2_2 _11354_ (.A(_05256_),
    .B(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hd__o32a_1 _11355_ (.A1(_05230_),
    .A2(_05243_),
    .A3(_05254_),
    .B1(_05255_),
    .B2(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__nor2_1 _11356_ (.A(_05242_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__xnor2_1 _11357_ (.A(_05242_),
    .B(_05260_),
    .Y(_05262_));
 sky130_fd_sc_hd__nor2_1 _11358_ (.A(_05258_),
    .B(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__nor3_1 _11359_ (.A(_05227_),
    .B(_05232_),
    .C(_05236_),
    .Y(_05264_));
 sky130_fd_sc_hd__nor2_1 _11360_ (.A(_05237_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__o21a_1 _11361_ (.A1(_05261_),
    .A2(_05263_),
    .B1(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__nor3_1 _11362_ (.A(_05261_),
    .B(_05263_),
    .C(_05265_),
    .Y(_05267_));
 sky130_fd_sc_hd__nor2_1 _11363_ (.A(_05266_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _11364_ (.A(_05258_),
    .B(_05262_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2b_1 _11365_ (.A_N(_05263_),
    .B(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__xor2_2 _11366_ (.A(_05255_),
    .B(_05259_),
    .X(_05271_));
 sky130_fd_sc_hd__xnor2_1 _11367_ (.A(_05250_),
    .B(_05252_),
    .Y(_05272_));
 sky130_fd_sc_hd__a22oi_1 _11368_ (.A1(net1471),
    .A2(net1668),
    .B1(net935),
    .B2(net1421),
    .Y(_05273_));
 sky130_fd_sc_hd__nor2_1 _11369_ (.A(_05253_),
    .B(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__and4_1 _11370_ (.A(net1421),
    .B(net1471),
    .C(net935),
    .D(net2132),
    .X(_05275_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(net1156),
    .B(net1668),
    .Y(_05276_));
 sky130_fd_sc_hd__a22o_1 _11372_ (.A1(net1471),
    .A2(net935),
    .B1(net2132),
    .B2(net1421),
    .X(_05277_));
 sky130_fd_sc_hd__and2b_1 _11373_ (.A_N(_05275_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__a31o_1 _11374_ (.A1(net1156),
    .A2(net1668),
    .A3(_05277_),
    .B1(_05275_),
    .X(_05279_));
 sky130_fd_sc_hd__a22oi_1 _11375_ (.A1(net1813),
    .A2(net1837),
    .B1(net2003),
    .B2(net1156),
    .Y(_05280_));
 sky130_fd_sc_hd__and4_1 _11376_ (.A(net1156),
    .B(net1813),
    .C(net1837),
    .D(net2003),
    .X(_05281_));
 sky130_fd_sc_hd__nor2_1 _11377_ (.A(_05280_),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hd__a21oi_1 _11378_ (.A1(net1995),
    .A2(net872),
    .B1(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__and3_1 _11379_ (.A(net1995),
    .B(net872),
    .C(_05282_),
    .X(_05284_));
 sky130_fd_sc_hd__or2_1 _11380_ (.A(_05283_),
    .B(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__xor2_2 _11381_ (.A(_05274_),
    .B(_05279_),
    .X(_05286_));
 sky130_fd_sc_hd__and2b_1 _11382_ (.A_N(_05285_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a21oi_1 _11383_ (.A1(_05274_),
    .A2(_05279_),
    .B1(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__o211a_1 _11384_ (.A1(_05281_),
    .A2(_05284_),
    .B1(net1995),
    .C1(net714),
    .X(_05289_));
 sky130_fd_sc_hd__a211oi_1 _11385_ (.A1(net1995),
    .A2(net714),
    .B1(_05281_),
    .C1(_05284_),
    .Y(_05290_));
 sky130_fd_sc_hd__or2_1 _11386_ (.A(_05289_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__xnor2_1 _11387_ (.A(_05272_),
    .B(_05288_),
    .Y(_05292_));
 sky130_fd_sc_hd__nor2_1 _11388_ (.A(_05291_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__o21ba_1 _11389_ (.A1(_05272_),
    .A2(_05288_),
    .B1_N(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__nand2b_1 _11390_ (.A_N(_05294_),
    .B(_05271_),
    .Y(_05295_));
 sky130_fd_sc_hd__xnor2_2 _11391_ (.A(_05271_),
    .B(_05294_),
    .Y(_05296_));
 sky130_fd_sc_hd__a21bo_1 _11392_ (.A1(_05289_),
    .A2(_05296_),
    .B1_N(_05295_),
    .X(_05297_));
 sky130_fd_sc_hd__and2b_1 _11393_ (.A_N(_05270_),
    .B(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__xor2_1 _11394_ (.A(_05270_),
    .B(_05297_),
    .X(_05299_));
 sky130_fd_sc_hd__inv_2 _11395_ (.A(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__xnor2_2 _11396_ (.A(_05289_),
    .B(_05296_),
    .Y(_05301_));
 sky130_fd_sc_hd__and2_1 _11397_ (.A(_05291_),
    .B(_05292_),
    .X(_05302_));
 sky130_fd_sc_hd__or2_1 _11398_ (.A(_05293_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__xor2_2 _11399_ (.A(_05285_),
    .B(_05286_),
    .X(_05304_));
 sky130_fd_sc_hd__xnor2_2 _11400_ (.A(_05276_),
    .B(_05278_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand4_1 _11401_ (.A(net1471),
    .B(net1156),
    .C(net935),
    .D(net2132),
    .Y(_05306_));
 sky130_fd_sc_hd__a22o_1 _11402_ (.A1(net1156),
    .A2(net935),
    .B1(net2132),
    .B2(net1471),
    .X(_05307_));
 sky130_fd_sc_hd__nand4_1 _11403_ (.A(net1995),
    .B(net1668),
    .C(_05306_),
    .D(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__and2_1 _11404_ (.A(_05306_),
    .B(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__nand2b_1 _11405_ (.A_N(_05309_),
    .B(_05305_),
    .Y(_05310_));
 sky130_fd_sc_hd__and4_1 _11406_ (.A(net1995),
    .B(net1721),
    .C(net1837),
    .D(net2003),
    .X(_05311_));
 sky130_fd_sc_hd__a22o_1 _11407_ (.A1(net1721),
    .A2(net1837),
    .B1(net2003),
    .B2(net1995),
    .X(_05312_));
 sky130_fd_sc_hd__inv_2 _11408_ (.A(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__and4b_1 _11409_ (.A_N(_05311_),
    .B(_05312_),
    .C(net2243),
    .D(net872),
    .X(_05314_));
 sky130_fd_sc_hd__o2bb2a_1 _11410_ (.A1_N(net2243),
    .A2_N(net872),
    .B1(_05311_),
    .B2(_05313_),
    .X(_05315_));
 sky130_fd_sc_hd__or2_1 _11411_ (.A(_05314_),
    .B(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__xnor2_2 _11412_ (.A(_05305_),
    .B(_05309_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand2b_1 _11413_ (.A_N(_05316_),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _11414_ (.A(_05310_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__a21oi_1 _11415_ (.A1(_05310_),
    .A2(_05318_),
    .B1(_05304_),
    .Y(_05320_));
 sky130_fd_sc_hd__o211a_1 _11416_ (.A1(_05311_),
    .A2(_05314_),
    .B1(net2243),
    .C1(net1741),
    .X(_05321_));
 sky130_fd_sc_hd__a211oi_1 _11417_ (.A1(net2243),
    .A2(net714),
    .B1(_05311_),
    .C1(_05314_),
    .Y(_05322_));
 sky130_fd_sc_hd__or2_1 _11418_ (.A(_05321_),
    .B(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__xnor2_2 _11419_ (.A(_05304_),
    .B(_05319_),
    .Y(_05324_));
 sky130_fd_sc_hd__and2b_1 _11420_ (.A_N(_05323_),
    .B(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__nor2_1 _11421_ (.A(_05320_),
    .B(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(_05303_),
    .B(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__xor2_2 _11423_ (.A(_05303_),
    .B(_05326_),
    .X(_05328_));
 sky130_fd_sc_hd__nand2_1 _11424_ (.A(_05321_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand2_1 _11425_ (.A(_05327_),
    .B(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2b_1 _11426_ (.A_N(_05330_),
    .B(_05301_),
    .Y(_05331_));
 sky130_fd_sc_hd__a21oi_1 _11427_ (.A1(_05327_),
    .A2(_05329_),
    .B1(_05301_),
    .Y(_05332_));
 sky130_fd_sc_hd__xnor2_2 _11428_ (.A(_05321_),
    .B(_05328_),
    .Y(_05333_));
 sky130_fd_sc_hd__xnor2_2 _11429_ (.A(_05323_),
    .B(_05324_),
    .Y(_05334_));
 sky130_fd_sc_hd__xnor2_2 _11430_ (.A(_05316_),
    .B(_05317_),
    .Y(_05335_));
 sky130_fd_sc_hd__a22o_1 _11431_ (.A1(net1995),
    .A2(net1668),
    .B1(_05306_),
    .B2(_05307_),
    .X(_05336_));
 sky130_fd_sc_hd__nand4_1 _11432_ (.A(net1156),
    .B(net1995),
    .C(net2361),
    .D(net2132),
    .Y(_05337_));
 sky130_fd_sc_hd__and2_1 _11433_ (.A(net2243),
    .B(net1668),
    .X(_05338_));
 sky130_fd_sc_hd__a22o_1 _11434_ (.A1(net1995),
    .A2(net2361),
    .B1(net2132),
    .B2(net1156),
    .X(_05339_));
 sky130_fd_sc_hd__nand3_1 _11435_ (.A(_05337_),
    .B(_05338_),
    .C(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21bo_1 _11436_ (.A1(_05338_),
    .A2(_05339_),
    .B1_N(_05337_),
    .X(_05341_));
 sky130_fd_sc_hd__and3_1 _11437_ (.A(_05308_),
    .B(_05336_),
    .C(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__and4_1 _11438_ (.A(net2243),
    .B(net1611),
    .C(net1837),
    .D(net2003),
    .X(_05343_));
 sky130_fd_sc_hd__a22o_1 _11439_ (.A1(net1611),
    .A2(net1837),
    .B1(net2003),
    .B2(net2243),
    .X(_05344_));
 sky130_fd_sc_hd__and2b_1 _11440_ (.A_N(_05343_),
    .B(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(net1813),
    .B(net872),
    .Y(_05346_));
 sky130_fd_sc_hd__xnor2_1 _11442_ (.A(_05345_),
    .B(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__a21oi_1 _11443_ (.A1(_05308_),
    .A2(_05336_),
    .B1(_05341_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor3b_1 _11444_ (.A(_05342_),
    .B(_05348_),
    .C_N(_05347_),
    .Y(_05349_));
 sky130_fd_sc_hd__nor2_1 _11445_ (.A(_05342_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2b_1 _11446_ (.A_N(_05350_),
    .B(_05335_),
    .Y(_05351_));
 sky130_fd_sc_hd__a31oi_2 _11447_ (.A1(net1813),
    .A2(net872),
    .A3(_05344_),
    .B1(_05343_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _11448_ (.A(net1813),
    .B(net1743),
    .Y(_05353_));
 sky130_fd_sc_hd__nor2_1 _11449_ (.A(_05352_),
    .B(_05353_),
    .Y(_05354_));
 sky130_fd_sc_hd__xnor2_1 _11450_ (.A(_05352_),
    .B(_05353_),
    .Y(_05355_));
 sky130_fd_sc_hd__and2b_1 _11451_ (.A_N(_05335_),
    .B(_05350_),
    .X(_05356_));
 sky130_fd_sc_hd__xnor2_1 _11452_ (.A(_05335_),
    .B(_05350_),
    .Y(_05357_));
 sky130_fd_sc_hd__o21a_1 _11453_ (.A1(_05355_),
    .A2(_05356_),
    .B1(_05351_),
    .X(_05358_));
 sky130_fd_sc_hd__and2b_1 _11454_ (.A_N(_05358_),
    .B(_05334_),
    .X(_05359_));
 sky130_fd_sc_hd__xnor2_2 _11455_ (.A(_05334_),
    .B(_05358_),
    .Y(_05360_));
 sky130_fd_sc_hd__a21o_1 _11456_ (.A1(_05354_),
    .A2(_05360_),
    .B1(_05359_),
    .X(_05361_));
 sky130_fd_sc_hd__and2b_1 _11457_ (.A_N(_05333_),
    .B(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__xnor2_2 _11458_ (.A(_05354_),
    .B(_05360_),
    .Y(_05363_));
 sky130_fd_sc_hd__xnor2_1 _11459_ (.A(_05355_),
    .B(_05357_),
    .Y(_05364_));
 sky130_fd_sc_hd__o21ba_1 _11460_ (.A1(_05342_),
    .A2(_05348_),
    .B1_N(_05347_),
    .X(_05365_));
 sky130_fd_sc_hd__a21o_1 _11461_ (.A1(_05337_),
    .A2(_05339_),
    .B1(_05338_),
    .X(_05366_));
 sky130_fd_sc_hd__nand4_2 _11462_ (.A(net1995),
    .B(net2243),
    .C(net2361),
    .D(net2132),
    .Y(_05367_));
 sky130_fd_sc_hd__and2_1 _11463_ (.A(net1813),
    .B(net1668),
    .X(_05368_));
 sky130_fd_sc_hd__a22o_1 _11464_ (.A1(net2243),
    .A2(net2361),
    .B1(net2132),
    .B2(net1995),
    .X(_05369_));
 sky130_fd_sc_hd__nand3_1 _11465_ (.A(_05367_),
    .B(_05368_),
    .C(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__a21bo_1 _11466_ (.A1(_05368_),
    .A2(_05369_),
    .B1_N(_05367_),
    .X(_05371_));
 sky130_fd_sc_hd__nand3_1 _11467_ (.A(_05340_),
    .B(_05366_),
    .C(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__a22oi_1 _11468_ (.A1(net1721),
    .A2(net872),
    .B1(net2003),
    .B2(net1813),
    .Y(_05373_));
 sky130_fd_sc_hd__and4_1 _11469_ (.A(net1813),
    .B(net1721),
    .C(net2838),
    .D(net2003),
    .X(_05374_));
 sky130_fd_sc_hd__nor2_1 _11470_ (.A(_05373_),
    .B(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__a21o_1 _11471_ (.A1(_05340_),
    .A2(_05366_),
    .B1(_05371_),
    .X(_05376_));
 sky130_fd_sc_hd__nand3_1 _11472_ (.A(_05372_),
    .B(_05375_),
    .C(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__a21bo_1 _11473_ (.A1(_05375_),
    .A2(_05376_),
    .B1_N(_05372_),
    .X(_05378_));
 sky130_fd_sc_hd__nor3b_1 _11474_ (.A(_05349_),
    .B(_05365_),
    .C_N(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__a21o_1 _11475_ (.A1(net1721),
    .A2(net1743),
    .B1(_05374_),
    .X(_05380_));
 sky130_fd_sc_hd__nand2_1 _11476_ (.A(net1743),
    .B(_05374_),
    .Y(_05381_));
 sky130_fd_sc_hd__nand4_1 _11477_ (.A(net1421),
    .B(net2239),
    .C(_05380_),
    .D(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__a22o_1 _11478_ (.A1(net1421),
    .A2(net2239),
    .B1(_05380_),
    .B2(_05381_),
    .X(_05383_));
 sky130_fd_sc_hd__and2_1 _11479_ (.A(_05382_),
    .B(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__o21ba_1 _11480_ (.A1(_05349_),
    .A2(_05365_),
    .B1_N(_05378_),
    .X(_05385_));
 sky130_fd_sc_hd__nor3b_1 _11481_ (.A(_05379_),
    .B(_05385_),
    .C_N(_05384_),
    .Y(_05386_));
 sky130_fd_sc_hd__or2_1 _11482_ (.A(_05379_),
    .B(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__nand2_1 _11483_ (.A(_05364_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _11484_ (.A(_05381_),
    .B(_05382_),
    .Y(_05389_));
 sky130_fd_sc_hd__xor2_1 _11485_ (.A(_05364_),
    .B(_05387_),
    .X(_05390_));
 sky130_fd_sc_hd__a21bo_1 _11486_ (.A1(_05389_),
    .A2(_05390_),
    .B1_N(_05388_),
    .X(_05391_));
 sky130_fd_sc_hd__and2b_1 _11487_ (.A_N(_05363_),
    .B(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__xnor2_2 _11488_ (.A(_05363_),
    .B(_05391_),
    .Y(_05393_));
 sky130_fd_sc_hd__xnor2_1 _11489_ (.A(_05389_),
    .B(_05390_),
    .Y(_05394_));
 sky130_fd_sc_hd__o21ba_1 _11490_ (.A1(_05379_),
    .A2(_05385_),
    .B1_N(_05384_),
    .X(_05395_));
 sky130_fd_sc_hd__a21o_1 _11491_ (.A1(_05372_),
    .A2(_05376_),
    .B1(_05375_),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _11492_ (.A1(_05367_),
    .A2(_05369_),
    .B1(_05368_),
    .X(_05397_));
 sky130_fd_sc_hd__nand4_1 _11493_ (.A(net2243),
    .B(net1813),
    .C(net935),
    .D(net2132),
    .Y(_05398_));
 sky130_fd_sc_hd__and2_1 _11494_ (.A(net1721),
    .B(net1668),
    .X(_05399_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(net1813),
    .A2(net935),
    .B1(net2132),
    .B2(net2243),
    .X(_05400_));
 sky130_fd_sc_hd__nand3_1 _11496_ (.A(_05398_),
    .B(_05399_),
    .C(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__a21bo_1 _11497_ (.A1(_05399_),
    .A2(_05400_),
    .B1_N(_05398_),
    .X(_05402_));
 sky130_fd_sc_hd__nand3_1 _11498_ (.A(_05370_),
    .B(_05397_),
    .C(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a22oi_1 _11499_ (.A1(net1611),
    .A2(net872),
    .B1(net2003),
    .B2(net1721),
    .Y(_05404_));
 sky130_fd_sc_hd__and4_1 _11500_ (.A(net1721),
    .B(net1611),
    .C(net872),
    .D(net2003),
    .X(_05405_));
 sky130_fd_sc_hd__nor2_1 _11501_ (.A(_05404_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__a21o_1 _11502_ (.A1(_05370_),
    .A2(_05397_),
    .B1(_05402_),
    .X(_05407_));
 sky130_fd_sc_hd__nand3_1 _11503_ (.A(_05403_),
    .B(_05406_),
    .C(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__a21bo_1 _11504_ (.A1(_05406_),
    .A2(_05407_),
    .B1_N(_05403_),
    .X(_05409_));
 sky130_fd_sc_hd__nand3_2 _11505_ (.A(_05377_),
    .B(_05396_),
    .C(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _11506_ (.A(net1471),
    .B(net2239),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _11507_ (.A(net1611),
    .B(net1743),
    .Y(_05412_));
 sky130_fd_sc_hd__mux2_1 _11508_ (.A0(_05412_),
    .A1(net1743),
    .S(_05405_),
    .X(_05413_));
 sky130_fd_sc_hd__xor2_1 _11509_ (.A(_05411_),
    .B(_05413_),
    .X(_05414_));
 sky130_fd_sc_hd__a21o_1 _11510_ (.A1(_05377_),
    .A2(_05396_),
    .B1(_05409_),
    .X(_05415_));
 sky130_fd_sc_hd__and3_1 _11511_ (.A(_05410_),
    .B(_05414_),
    .C(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__nand3_1 _11512_ (.A(_05410_),
    .B(_05414_),
    .C(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__a211o_1 _11513_ (.A1(_05410_),
    .A2(_05417_),
    .B1(_05386_),
    .C1(_05395_),
    .X(_05418_));
 sky130_fd_sc_hd__o2bb2ai_1 _11514_ (.A1_N(net1743),
    .A2_N(_05405_),
    .B1(_05411_),
    .B2(_05413_),
    .Y(_05419_));
 sky130_fd_sc_hd__o211ai_1 _11515_ (.A1(_05386_),
    .A2(_05395_),
    .B1(_05410_),
    .C1(_05417_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand3_1 _11516_ (.A(_05418_),
    .B(_05419_),
    .C(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(_05418_),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__and2b_1 _11518_ (.A_N(_05394_),
    .B(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__xnor2_1 _11519_ (.A(_05394_),
    .B(_05422_),
    .Y(_05424_));
 sky130_fd_sc_hd__a21o_1 _11520_ (.A1(_05418_),
    .A2(_05420_),
    .B1(_05419_),
    .X(_05425_));
 sky130_fd_sc_hd__and2_1 _11521_ (.A(_05421_),
    .B(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__a21o_1 _11522_ (.A1(_05403_),
    .A2(_05407_),
    .B1(_05406_),
    .X(_05427_));
 sky130_fd_sc_hd__a21o_1 _11523_ (.A1(_05398_),
    .A2(_05400_),
    .B1(_05399_),
    .X(_05428_));
 sky130_fd_sc_hd__and3_1 _11524_ (.A(net1813),
    .B(net1721),
    .C(net2132),
    .X(_05429_));
 sky130_fd_sc_hd__nand2_1 _11525_ (.A(net1611),
    .B(net1668),
    .Y(_05430_));
 sky130_fd_sc_hd__a22o_1 _11526_ (.A1(net1721),
    .A2(net935),
    .B1(net2132),
    .B2(net1813),
    .X(_05431_));
 sky130_fd_sc_hd__a21bo_1 _11527_ (.A1(net935),
    .A2(_05429_),
    .B1_N(_05431_),
    .X(_05432_));
 sky130_fd_sc_hd__a32o_1 _11528_ (.A1(net1611),
    .A2(net1668),
    .A3(_05431_),
    .B1(_05429_),
    .B2(net935),
    .X(_05433_));
 sky130_fd_sc_hd__nand3_1 _11529_ (.A(_05401_),
    .B(_05428_),
    .C(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(net1611),
    .B(net2003),
    .X(_05435_));
 sky130_fd_sc_hd__a21o_1 _11531_ (.A1(_05401_),
    .A2(_05428_),
    .B1(_05433_),
    .X(_05436_));
 sky130_fd_sc_hd__nand3_1 _11532_ (.A(_05434_),
    .B(_05435_),
    .C(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21bo_1 _11533_ (.A1(_05435_),
    .A2(_05436_),
    .B1_N(_05434_),
    .X(_05438_));
 sky130_fd_sc_hd__nand3_2 _11534_ (.A(_05408_),
    .B(_05427_),
    .C(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__a21o_1 _11535_ (.A1(_05408_),
    .A2(_05427_),
    .B1(_05438_),
    .X(_05440_));
 sky130_fd_sc_hd__nand4_2 _11536_ (.A(net1156),
    .B(net2239),
    .C(_05439_),
    .D(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__a21oi_1 _11537_ (.A1(_05410_),
    .A2(_05415_),
    .B1(_05414_),
    .Y(_05442_));
 sky130_fd_sc_hd__a211o_1 _11538_ (.A1(_05439_),
    .A2(_05441_),
    .B1(_05442_),
    .C1(_05416_),
    .X(_05443_));
 sky130_fd_sc_hd__inv_2 _11539_ (.A(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__a22o_1 _11540_ (.A1(net1156),
    .A2(net2239),
    .B1(_05439_),
    .B2(_05440_),
    .X(_05445_));
 sky130_fd_sc_hd__a21o_1 _11541_ (.A1(_05434_),
    .A2(_05436_),
    .B1(_05435_),
    .X(_05446_));
 sky130_fd_sc_hd__xor2_2 _11542_ (.A(_05430_),
    .B(_05432_),
    .X(_05447_));
 sky130_fd_sc_hd__and3_1 _11543_ (.A(net1721),
    .B(net1611),
    .C(net2132),
    .X(_05448_));
 sky130_fd_sc_hd__nand2_2 _11544_ (.A(net935),
    .B(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__and3_1 _11545_ (.A(net935),
    .B(_05447_),
    .C(_05448_),
    .X(_05450_));
 sky130_fd_sc_hd__nand3_1 _11546_ (.A(_05437_),
    .B(_05446_),
    .C(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__and2_1 _11547_ (.A(net1995),
    .B(net2239),
    .X(_05452_));
 sky130_fd_sc_hd__a21o_1 _11548_ (.A1(_05437_),
    .A2(_05446_),
    .B1(_05450_),
    .X(_05453_));
 sky130_fd_sc_hd__nand3_1 _11549_ (.A(_05451_),
    .B(_05452_),
    .C(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21bo_1 _11550_ (.A1(_05452_),
    .A2(_05453_),
    .B1_N(_05451_),
    .X(_05455_));
 sky130_fd_sc_hd__and3_1 _11551_ (.A(_05441_),
    .B(_05445_),
    .C(_05455_),
    .X(_05456_));
 sky130_fd_sc_hd__o211ai_1 _11552_ (.A1(_05416_),
    .A2(_05442_),
    .B1(_05441_),
    .C1(_05439_),
    .Y(_05457_));
 sky130_fd_sc_hd__and3_1 _11553_ (.A(_05443_),
    .B(_05456_),
    .C(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__or2_1 _11554_ (.A(_05444_),
    .B(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__a21o_1 _11555_ (.A1(_05421_),
    .A2(_05425_),
    .B1(_05444_),
    .X(_05460_));
 sky130_fd_sc_hd__a21oi_1 _11556_ (.A1(_05443_),
    .A2(_05457_),
    .B1(_05456_),
    .Y(_05461_));
 sky130_fd_sc_hd__nor2_2 _11557_ (.A(_05458_),
    .B(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__a21o_1 _11558_ (.A1(_05451_),
    .A2(_05453_),
    .B1(_05452_),
    .X(_05463_));
 sky130_fd_sc_hd__and2_1 _11559_ (.A(_05454_),
    .B(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__xnor2_2 _11560_ (.A(_05447_),
    .B(_05449_),
    .Y(_05465_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(net2243),
    .B(net2239),
    .Y(_05466_));
 sky130_fd_sc_hd__and3_1 _11562_ (.A(net2243),
    .B(net2239),
    .C(_05465_),
    .X(_05467_));
 sky130_fd_sc_hd__a21oi_1 _11563_ (.A1(_05441_),
    .A2(_05445_),
    .B1(_05455_),
    .Y(_05468_));
 sky130_fd_sc_hd__a2bb2o_1 _11564_ (.A1_N(_05456_),
    .A2_N(_05468_),
    .B1(_05467_),
    .B2(_05464_),
    .X(_05469_));
 sky130_fd_sc_hd__inv_2 _11565_ (.A(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__and4bb_1 _11566_ (.A_N(_05456_),
    .B_N(_05468_),
    .C(_05467_),
    .D(_05464_),
    .X(_05471_));
 sky130_fd_sc_hd__xor2_2 _11567_ (.A(_05465_),
    .B(_05466_),
    .X(_05472_));
 sky130_fd_sc_hd__a22o_1 _11568_ (.A1(net1611),
    .A2(net935),
    .B1(net2132),
    .B2(net1721),
    .X(_05473_));
 sky130_fd_sc_hd__nand4_2 _11569_ (.A(net1813),
    .B(net2239),
    .C(_05449_),
    .D(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a22o_1 _11570_ (.A1(net1813),
    .A2(net2239),
    .B1(_05449_),
    .B2(_05473_),
    .X(_05475_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(_05474_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__and2_1 _11572_ (.A(net2239),
    .B(_05448_),
    .X(_05477_));
 sky130_fd_sc_hd__and4b_1 _11573_ (.A_N(_05472_),
    .B(_05474_),
    .C(_05475_),
    .D(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__inv_2 _11574_ (.A(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__o21bai_1 _11575_ (.A1(_05472_),
    .A2(_05474_),
    .B1_N(_05467_),
    .Y(_05480_));
 sky130_fd_sc_hd__and3_1 _11576_ (.A(_05454_),
    .B(_05463_),
    .C(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _11577_ (.A1(_05454_),
    .A2(_05463_),
    .B1(_05480_),
    .Y(_05482_));
 sky130_fd_sc_hd__nor2_1 _11578_ (.A(_05481_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__or4bb_1 _11579_ (.A(_05472_),
    .B(_05474_),
    .C_N(_05454_),
    .D_N(_05463_),
    .X(_05484_));
 sky130_fd_sc_hd__o31ai_2 _11580_ (.A1(_05479_),
    .A2(_05481_),
    .A3(_05482_),
    .B1(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__o21a_1 _11581_ (.A1(_05471_),
    .A2(_05485_),
    .B1(_05469_),
    .X(_05486_));
 sky130_fd_sc_hd__a32o_1 _11582_ (.A1(_05460_),
    .A2(_05462_),
    .A3(_05486_),
    .B1(_05459_),
    .B2(_05426_),
    .X(_05487_));
 sky130_fd_sc_hd__a21o_1 _11583_ (.A1(_05424_),
    .A2(_05487_),
    .B1(_05423_),
    .X(_05488_));
 sky130_fd_sc_hd__a21o_2 _11584_ (.A1(_05393_),
    .A2(_05488_),
    .B1(_05392_),
    .X(_05489_));
 sky130_fd_sc_hd__xnor2_2 _11585_ (.A(_05333_),
    .B(_05361_),
    .Y(_05490_));
 sky130_fd_sc_hd__a21o_1 _11586_ (.A1(_05489_),
    .A2(_05490_),
    .B1(_05362_),
    .X(_05491_));
 sky130_fd_sc_hd__a211o_1 _11587_ (.A1(_05489_),
    .A2(_05490_),
    .B1(_05332_),
    .C1(_05362_),
    .X(_05492_));
 sky130_fd_sc_hd__and3_1 _11588_ (.A(_05300_),
    .B(_05331_),
    .C(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__a31o_1 _11589_ (.A1(_05300_),
    .A2(_05331_),
    .A3(_05492_),
    .B1(_05298_),
    .X(_05494_));
 sky130_fd_sc_hd__a21oi_2 _11590_ (.A1(_05268_),
    .A2(_05494_),
    .B1(_05266_),
    .Y(_05495_));
 sky130_fd_sc_hd__nor2_1 _11591_ (.A(_05240_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__xnor2_2 _11592_ (.A(_05240_),
    .B(_05495_),
    .Y(_05497_));
 sky130_fd_sc_hd__xor2_2 _11593_ (.A(_05220_),
    .B(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__xor2_2 _11594_ (.A(_04701_),
    .B(_04936_),
    .X(_05499_));
 sky130_fd_sc_hd__xor2_4 _11595_ (.A(_05003_),
    .B(_05215_),
    .X(_05500_));
 sky130_fd_sc_hd__xnor2_1 _11596_ (.A(_05268_),
    .B(_05494_),
    .Y(_05501_));
 sky130_fd_sc_hd__xnor2_1 _11597_ (.A(_05499_),
    .B(_05500_),
    .Y(_05502_));
 sky130_fd_sc_hd__nor2_1 _11598_ (.A(_05501_),
    .B(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__a21oi_2 _11599_ (.A1(_05499_),
    .A2(_05500_),
    .B1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2b_1 _11600_ (.A_N(_05504_),
    .B(_05498_),
    .Y(_05505_));
 sky130_fd_sc_hd__xnor2_2 _11601_ (.A(_05498_),
    .B(_05504_),
    .Y(_05506_));
 sky130_fd_sc_hd__nand3_1 _11602_ (.A(_04656_),
    .B(_04657_),
    .C(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__a21o_1 _11603_ (.A1(_04656_),
    .A2(_04657_),
    .B1(_05506_),
    .X(_05508_));
 sky130_fd_sc_hd__and2_1 _11604_ (.A(_05501_),
    .B(_05502_),
    .X(_05509_));
 sky130_fd_sc_hd__or2_1 _11605_ (.A(_05503_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__a21oi_1 _11606_ (.A1(_04766_),
    .A2(_04934_),
    .B1(_04732_),
    .Y(_05511_));
 sky130_fd_sc_hd__xnor2_2 _11607_ (.A(_05029_),
    .B(_05214_),
    .Y(_05512_));
 sky130_fd_sc_hd__or3_1 _11608_ (.A(_04935_),
    .B(_05511_),
    .C(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__a21oi_1 _11609_ (.A1(_05331_),
    .A2(_05492_),
    .B1(_05300_),
    .Y(_05514_));
 sky130_fd_sc_hd__nor2_2 _11610_ (.A(_05493_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_1 _11611_ (.A1(_04935_),
    .A2(_05511_),
    .B1(_05512_),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_1 _11612_ (.A(_05513_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__a21bo_1 _11613_ (.A1(_05515_),
    .A2(_05516_),
    .B1_N(_05513_),
    .X(_05518_));
 sky130_fd_sc_hd__and2b_1 _11614_ (.A_N(_05510_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__a22oi_1 _11615_ (.A1(_04617_),
    .A2(_04618_),
    .B1(_04619_),
    .B2(_04605_),
    .Y(_05520_));
 sky130_fd_sc_hd__nor2_1 _11616_ (.A(_04620_),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__xor2_2 _11617_ (.A(_05510_),
    .B(_05518_),
    .X(_05522_));
 sky130_fd_sc_hd__nor3_1 _11618_ (.A(_04620_),
    .B(_05520_),
    .C(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__o211a_1 _11619_ (.A1(_05519_),
    .A2(_05523_),
    .B1(_05507_),
    .C1(_05508_),
    .X(_05524_));
 sky130_fd_sc_hd__a211oi_1 _11620_ (.A1(_05507_),
    .A2(_05508_),
    .B1(_05519_),
    .C1(_05523_),
    .Y(_05525_));
 sky130_fd_sc_hd__nor3_1 _11621_ (.A(_04632_),
    .B(_05524_),
    .C(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21a_1 _11622_ (.A1(_05524_),
    .A2(_05525_),
    .B1(_04632_),
    .X(_05527_));
 sky130_fd_sc_hd__xnor2_1 _11623_ (.A(_05521_),
    .B(_05522_),
    .Y(_05528_));
 sky130_fd_sc_hd__xnor2_2 _11624_ (.A(_05515_),
    .B(_05517_),
    .Y(_05529_));
 sky130_fd_sc_hd__a31o_1 _11625_ (.A1(_05085_),
    .A2(_05112_),
    .A3(_05212_),
    .B1(_05081_),
    .X(_05530_));
 sky130_fd_sc_hd__or2_1 _11626_ (.A(_05030_),
    .B(_05052_),
    .X(_05531_));
 sky130_fd_sc_hd__and2_1 _11627_ (.A(_05084_),
    .B(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__xnor2_2 _11628_ (.A(_05530_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__and2_1 _11629_ (.A(_04766_),
    .B(_04768_),
    .X(_05534_));
 sky130_fd_sc_hd__xnor2_2 _11630_ (.A(_04933_),
    .B(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__or2_1 _11631_ (.A(_05533_),
    .B(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__xnor2_2 _11632_ (.A(_05533_),
    .B(_05535_),
    .Y(_05537_));
 sky130_fd_sc_hd__xnor2_1 _11633_ (.A(_05301_),
    .B(_05330_),
    .Y(_05538_));
 sky130_fd_sc_hd__xnor2_2 _11634_ (.A(_05491_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__o21a_1 _11635_ (.A1(_05537_),
    .A2(_05539_),
    .B1(_05536_),
    .X(_05540_));
 sky130_fd_sc_hd__nand2b_1 _11636_ (.A_N(_05540_),
    .B(_05529_),
    .Y(_05541_));
 sky130_fd_sc_hd__xor2_1 _11637_ (.A(_04032_),
    .B(_04033_),
    .X(_05542_));
 sky130_fd_sc_hd__xnor2_2 _11638_ (.A(_05529_),
    .B(_05540_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand2_1 _11639_ (.A(_05542_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__a21bo_1 _11640_ (.A1(_05541_),
    .A2(_05544_),
    .B1_N(_05528_),
    .X(_05545_));
 sky130_fd_sc_hd__xor2_1 _11641_ (.A(_04568_),
    .B(_04570_),
    .X(_05546_));
 sky130_fd_sc_hd__nand3b_1 _11642_ (.A_N(_05528_),
    .B(_05541_),
    .C(_05544_),
    .Y(_05547_));
 sky130_fd_sc_hd__and3_1 _11643_ (.A(_05545_),
    .B(_05546_),
    .C(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__nand3_1 _11644_ (.A(_05545_),
    .B(_05546_),
    .C(_05547_),
    .Y(_05549_));
 sky130_fd_sc_hd__a211oi_1 _11645_ (.A1(_05545_),
    .A2(_05549_),
    .B1(_05526_),
    .C1(_05527_),
    .Y(_05550_));
 sky130_fd_sc_hd__o211a_1 _11646_ (.A1(_05526_),
    .A2(_05527_),
    .B1(_05545_),
    .C1(_05549_),
    .X(_05551_));
 sky130_fd_sc_hd__nor2_1 _11647_ (.A(_05550_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__xnor2_1 _11648_ (.A(_04571_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__a21oi_1 _11649_ (.A1(_05545_),
    .A2(_05547_),
    .B1(_05546_),
    .Y(_05554_));
 sky130_fd_sc_hd__xor2_1 _11650_ (.A(_05542_),
    .B(_05543_),
    .X(_05555_));
 sky130_fd_sc_hd__xnor2_2 _11651_ (.A(_05537_),
    .B(_05539_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21oi_2 _11652_ (.A1(_04827_),
    .A2(_04931_),
    .B1(_04798_),
    .Y(_05557_));
 sky130_fd_sc_hd__a21oi_2 _11653_ (.A1(_05112_),
    .A2(_05212_),
    .B1(_05085_),
    .Y(_05558_));
 sky130_fd_sc_hd__or4_2 _11654_ (.A(_04932_),
    .B(_05213_),
    .C(_05557_),
    .D(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__xor2_2 _11655_ (.A(_05489_),
    .B(_05490_),
    .X(_05560_));
 sky130_fd_sc_hd__o22ai_4 _11656_ (.A1(_04932_),
    .A2(_05557_),
    .B1(_05558_),
    .B2(_05213_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand3_1 _11657_ (.A(_05559_),
    .B(_05560_),
    .C(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _11658_ (.A(_05559_),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2b_1 _11659_ (.A_N(_05556_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(_03365_),
    .B(_03366_),
    .Y(_05565_));
 sky130_fd_sc_hd__nand2_2 _11661_ (.A(_03367_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__xnor2_4 _11662_ (.A(_03524_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_03617_),
    .B(_03618_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_2 _11664_ (.A(_03619_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__xnor2_4 _11665_ (.A(_03777_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__or2_1 _11666_ (.A(_05567_),
    .B(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__xor2_2 _11667_ (.A(_05567_),
    .B(_05570_),
    .X(_05572_));
 sky130_fd_sc_hd__xnor2_1 _11668_ (.A(_03875_),
    .B(_04028_),
    .Y(_05573_));
 sky130_fd_sc_hd__xnor2_2 _11669_ (.A(_03874_),
    .B(_05573_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_05572_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__xnor2_2 _11671_ (.A(_05572_),
    .B(_05574_),
    .Y(_05576_));
 sky130_fd_sc_hd__xor2_2 _11672_ (.A(_05556_),
    .B(_05563_),
    .X(_05577_));
 sky130_fd_sc_hd__o21ai_1 _11673_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05564_),
    .Y(_05578_));
 sky130_fd_sc_hd__nand2_1 _11674_ (.A(_05555_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand3_1 _11675_ (.A(_04373_),
    .B(_04409_),
    .C(_04564_),
    .Y(_05580_));
 sky130_fd_sc_hd__nand2_2 _11676_ (.A(_04565_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__xnor2_2 _11677_ (.A(_04120_),
    .B(_04299_),
    .Y(_05582_));
 sky130_fd_sc_hd__a21o_1 _11678_ (.A1(_05571_),
    .A2(_05575_),
    .B1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__nand3_1 _11679_ (.A(_05571_),
    .B(_05575_),
    .C(_05582_),
    .Y(_05584_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(_05583_),
    .B(_05584_),
    .Y(_05585_));
 sky130_fd_sc_hd__or2_1 _11681_ (.A(_05581_),
    .B(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__and2_1 _11682_ (.A(_05581_),
    .B(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__xor2_1 _11683_ (.A(_05581_),
    .B(_05585_),
    .X(_05588_));
 sky130_fd_sc_hd__xnor2_1 _11684_ (.A(_05555_),
    .B(_05578_),
    .Y(_05589_));
 sky130_fd_sc_hd__or3b_1 _11685_ (.A(_05589_),
    .B(_05587_),
    .C_N(_05586_),
    .X(_05590_));
 sky130_fd_sc_hd__a211oi_2 _11686_ (.A1(_05579_),
    .A2(_05590_),
    .B1(_05548_),
    .C1(_05554_),
    .Y(_05591_));
 sky130_fd_sc_hd__o211a_1 _11687_ (.A1(_05548_),
    .A2(_05554_),
    .B1(net3716),
    .C1(_05590_),
    .X(_05592_));
 sky130_fd_sc_hd__a211oi_2 _11688_ (.A1(net3686),
    .A2(_05586_),
    .B1(_05591_),
    .C1(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__or2_1 _11689_ (.A(_05591_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__and2b_1 _11690_ (.A_N(_05553_),
    .B(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__xnor2_1 _11691_ (.A(_05553_),
    .B(_05594_),
    .Y(_05596_));
 sky130_fd_sc_hd__o211a_1 _11692_ (.A1(_05591_),
    .A2(_05592_),
    .B1(net3686),
    .C1(_05586_),
    .X(_05597_));
 sky130_fd_sc_hd__xnor2_1 _11693_ (.A(_05588_),
    .B(_05589_),
    .Y(_05598_));
 sky130_fd_sc_hd__xnor2_2 _11694_ (.A(_05576_),
    .B(_05577_),
    .Y(_05599_));
 sky130_fd_sc_hd__a21o_1 _11695_ (.A1(_05559_),
    .A2(_05561_),
    .B1(_05560_),
    .X(_05600_));
 sky130_fd_sc_hd__nor2_1 _11696_ (.A(_04826_),
    .B(_04828_),
    .Y(_05601_));
 sky130_fd_sc_hd__xnor2_2 _11697_ (.A(_04930_),
    .B(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__or2_1 _11698_ (.A(_05111_),
    .B(_05113_),
    .X(_05603_));
 sky130_fd_sc_hd__xnor2_2 _11699_ (.A(_05211_),
    .B(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__and2_1 _11700_ (.A(_05602_),
    .B(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__xnor2_2 _11701_ (.A(_05393_),
    .B(_05488_),
    .Y(_05606_));
 sky130_fd_sc_hd__xnor2_2 _11702_ (.A(_05602_),
    .B(_05604_),
    .Y(_05607_));
 sky130_fd_sc_hd__nor2_1 _11703_ (.A(_05606_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__o211ai_2 _11704_ (.A1(_05605_),
    .A2(_05608_),
    .B1(_05562_),
    .C1(_05600_),
    .Y(_05609_));
 sky130_fd_sc_hd__xnor2_2 _11705_ (.A(_03903_),
    .B(_04027_),
    .Y(_05610_));
 sky130_fd_sc_hd__xor2_2 _11706_ (.A(_03521_),
    .B(_03523_),
    .X(_05611_));
 sky130_fd_sc_hd__xnor2_2 _11707_ (.A(_03774_),
    .B(_03776_),
    .Y(_05612_));
 sky130_fd_sc_hd__and2_1 _11708_ (.A(_05611_),
    .B(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__xnor2_1 _11709_ (.A(_05611_),
    .B(_05612_),
    .Y(_05614_));
 sky130_fd_sc_hd__nor2_1 _11710_ (.A(_05610_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__xor2_1 _11711_ (.A(_05610_),
    .B(_05614_),
    .X(_05616_));
 sky130_fd_sc_hd__a211o_1 _11712_ (.A1(_05562_),
    .A2(_05600_),
    .B1(_05605_),
    .C1(_05608_),
    .X(_05617_));
 sky130_fd_sc_hd__nand3_1 _11713_ (.A(_05609_),
    .B(_05616_),
    .C(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__and2_1 _11714_ (.A(_05609_),
    .B(_05618_),
    .X(_05619_));
 sky130_fd_sc_hd__or2_1 _11715_ (.A(_05599_),
    .B(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__or3_1 _11716_ (.A(_04411_),
    .B(_04445_),
    .C(_04563_),
    .X(_05621_));
 sky130_fd_sc_hd__and2_2 _11717_ (.A(_04564_),
    .B(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__nor3_1 _11718_ (.A(_04143_),
    .B(_04170_),
    .C(_04297_),
    .Y(_05623_));
 sky130_fd_sc_hd__nor2_1 _11719_ (.A(_04298_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21a_1 _11720_ (.A1(_05613_),
    .A2(_05615_),
    .B1(_05624_),
    .X(_05625_));
 sky130_fd_sc_hd__nor3_1 _11721_ (.A(_05613_),
    .B(_05615_),
    .C(_05624_),
    .Y(_05626_));
 sky130_fd_sc_hd__nor2_1 _11722_ (.A(_05625_),
    .B(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__xnor2_2 _11723_ (.A(_05622_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__xnor2_2 _11724_ (.A(_05599_),
    .B(_05619_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21a_1 _11725_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_05620_),
    .X(_05630_));
 sky130_fd_sc_hd__nand2b_1 _11726_ (.A_N(_05630_),
    .B(_05598_),
    .Y(_05631_));
 sky130_fd_sc_hd__a21o_1 _11727_ (.A1(_05622_),
    .A2(_05627_),
    .B1(net3799),
    .X(_05632_));
 sky130_fd_sc_hd__xnor2_1 _11728_ (.A(_05598_),
    .B(_05630_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_1 _11729_ (.A(_05632_),
    .B(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__o211a_1 _11730_ (.A1(_05593_),
    .A2(_05597_),
    .B1(_05631_),
    .C1(_05634_),
    .X(_05635_));
 sky130_fd_sc_hd__a211oi_1 _11731_ (.A1(_05631_),
    .A2(_05634_),
    .B1(_05593_),
    .C1(_05597_),
    .Y(_05636_));
 sky130_fd_sc_hd__xnor2_1 _11732_ (.A(_05632_),
    .B(_05633_),
    .Y(_05637_));
 sky130_fd_sc_hd__xor2_2 _11733_ (.A(_05628_),
    .B(_05629_),
    .X(_05638_));
 sky130_fd_sc_hd__a21o_1 _11734_ (.A1(_05609_),
    .A2(_05617_),
    .B1(_05616_),
    .X(_05639_));
 sky130_fd_sc_hd__xor2_2 _11735_ (.A(_05606_),
    .B(_05607_),
    .X(_05640_));
 sky130_fd_sc_hd__xor2_2 _11736_ (.A(net3214),
    .B(_04929_),
    .X(_05641_));
 sky130_fd_sc_hd__xor2_4 _11737_ (.A(_05209_),
    .B(_05210_),
    .X(_05642_));
 sky130_fd_sc_hd__xor2_1 _11738_ (.A(_05424_),
    .B(_05487_),
    .X(_05643_));
 sky130_fd_sc_hd__xor2_1 _11739_ (.A(net3215),
    .B(_05642_),
    .X(_05644_));
 sky130_fd_sc_hd__and2_1 _11740_ (.A(_05643_),
    .B(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__a21oi_2 _11741_ (.A1(_05641_),
    .A2(_05642_),
    .B1(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__and2b_1 _11742_ (.A_N(_05646_),
    .B(_05640_),
    .X(_05647_));
 sky130_fd_sc_hd__xnor2_2 _11743_ (.A(_03930_),
    .B(_04026_),
    .Y(_05648_));
 sky130_fd_sc_hd__xnor2_4 _11744_ (.A(_03423_),
    .B(_03520_),
    .Y(_05649_));
 sky130_fd_sc_hd__xor2_4 _11745_ (.A(_03677_),
    .B(_03773_),
    .X(_05650_));
 sky130_fd_sc_hd__xor2_2 _11746_ (.A(_05649_),
    .B(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2b_1 _11747_ (.A_N(_05648_),
    .B(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__xnor2_2 _11748_ (.A(_05648_),
    .B(_05651_),
    .Y(_05653_));
 sky130_fd_sc_hd__xnor2_2 _11749_ (.A(_05640_),
    .B(_05646_),
    .Y(_05654_));
 sky130_fd_sc_hd__and2_1 _11750_ (.A(_05653_),
    .B(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__o211ai_2 _11751_ (.A1(_05647_),
    .A2(_05655_),
    .B1(_05618_),
    .C1(_05639_),
    .Y(_05656_));
 sky130_fd_sc_hd__nor3_1 _11752_ (.A(_04446_),
    .B(_04477_),
    .C(_04562_),
    .Y(_05657_));
 sky130_fd_sc_hd__nor2_1 _11753_ (.A(_04563_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_2 _11754_ (.A1(_05649_),
    .A2(_05650_),
    .B1(_05652_),
    .Y(_05659_));
 sky130_fd_sc_hd__and3_1 _11755_ (.A(_04172_),
    .B(_04199_),
    .C(_04296_),
    .X(_05660_));
 sky130_fd_sc_hd__or2_1 _11756_ (.A(_04297_),
    .B(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__and2b_1 _11757_ (.A_N(_05661_),
    .B(_05659_),
    .X(_05662_));
 sky130_fd_sc_hd__xnor2_1 _11758_ (.A(_05659_),
    .B(_05661_),
    .Y(_05663_));
 sky130_fd_sc_hd__xor2_1 _11759_ (.A(_05658_),
    .B(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__a211o_1 _11760_ (.A1(_05618_),
    .A2(_05639_),
    .B1(_05647_),
    .C1(_05655_),
    .X(_05665_));
 sky130_fd_sc_hd__and3_1 _11761_ (.A(_05656_),
    .B(_05664_),
    .C(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a21boi_2 _11762_ (.A1(_05664_),
    .A2(_05665_),
    .B1_N(_05656_),
    .Y(_05667_));
 sky130_fd_sc_hd__and2b_1 _11763_ (.A_N(_05667_),
    .B(_05638_),
    .X(_05668_));
 sky130_fd_sc_hd__a21o_1 _11764_ (.A1(_05658_),
    .A2(_05663_),
    .B1(_05662_),
    .X(_05669_));
 sky130_fd_sc_hd__xnor2_2 _11765_ (.A(_05638_),
    .B(_05667_),
    .Y(_05670_));
 sky130_fd_sc_hd__a21oi_1 _11766_ (.A1(_05669_),
    .A2(_05670_),
    .B1(_05668_),
    .Y(_05671_));
 sky130_fd_sc_hd__or2_1 _11767_ (.A(_05637_),
    .B(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__xnor2_2 _11768_ (.A(_05669_),
    .B(_05670_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21oi_1 _11769_ (.A1(_05656_),
    .A2(_05665_),
    .B1(_05664_),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_1 _11770_ (.A(_05666_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__xnor2_2 _11771_ (.A(_05653_),
    .B(_05654_),
    .Y(_05676_));
 sky130_fd_sc_hd__nor2_1 _11772_ (.A(_03956_),
    .B(_04024_),
    .Y(_05677_));
 sky130_fd_sc_hd__nor2_1 _11773_ (.A(_04025_),
    .B(_05677_),
    .Y(_05678_));
 sky130_fd_sc_hd__xor2_2 _11774_ (.A(_03450_),
    .B(_03519_),
    .X(_05679_));
 sky130_fd_sc_hd__xor2_2 _11775_ (.A(_03704_),
    .B(_03772_),
    .X(_05680_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_05679_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__or2_1 _11777_ (.A(_05679_),
    .B(_05680_),
    .X(_05682_));
 sky130_fd_sc_hd__nand2_1 _11778_ (.A(_05681_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__xor2_2 _11779_ (.A(_05678_),
    .B(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__nor2_1 _11780_ (.A(_05643_),
    .B(_05644_),
    .Y(_05685_));
 sky130_fd_sc_hd__or2_2 _11781_ (.A(_05645_),
    .B(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__nor2_1 _11782_ (.A(_05684_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__and3_1 _11783_ (.A(_04479_),
    .B(_04505_),
    .C(_04561_),
    .X(_05688_));
 sky130_fd_sc_hd__nor2_1 _11784_ (.A(_04562_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__o31ai_2 _11785_ (.A1(_04025_),
    .A2(_05677_),
    .A3(_05683_),
    .B1(_05681_),
    .Y(_05690_));
 sky130_fd_sc_hd__or3_1 _11786_ (.A(_04200_),
    .B(_04225_),
    .C(_04295_),
    .X(_05691_));
 sky130_fd_sc_hd__nand2_1 _11787_ (.A(_04296_),
    .B(_05691_),
    .Y(_05692_));
 sky130_fd_sc_hd__and3_1 _11788_ (.A(_04296_),
    .B(_05690_),
    .C(_05691_),
    .X(_05693_));
 sky130_fd_sc_hd__xnor2_1 _11789_ (.A(_05690_),
    .B(_05692_),
    .Y(_05694_));
 sky130_fd_sc_hd__xor2_1 _11790_ (.A(_05689_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__xnor2_1 _11791_ (.A(_05676_),
    .B(_05687_),
    .Y(_05696_));
 sky130_fd_sc_hd__nand2_1 _11792_ (.A(_05695_),
    .B(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__o31ai_2 _11793_ (.A1(_05676_),
    .A2(_05684_),
    .A3(_05686_),
    .B1(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(_05675_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__a21oi_1 _11795_ (.A1(_05689_),
    .A2(_05694_),
    .B1(_05693_),
    .Y(_05700_));
 sky130_fd_sc_hd__xnor2_1 _11796_ (.A(_05675_),
    .B(_05698_),
    .Y(_05701_));
 sky130_fd_sc_hd__o21a_1 _11797_ (.A1(_05700_),
    .A2(_05701_),
    .B1(_05699_),
    .X(_05702_));
 sky130_fd_sc_hd__nor2_1 _11798_ (.A(_05673_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__xnor2_1 _11799_ (.A(_05700_),
    .B(_05701_),
    .Y(_05704_));
 sky130_fd_sc_hd__or2_1 _11800_ (.A(_05695_),
    .B(_05696_),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(_05697_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__o211a_1 _11802_ (.A1(_04225_),
    .A2(_04226_),
    .B1(_04247_),
    .C1(_04294_),
    .X(_05707_));
 sky130_fd_sc_hd__nor2_1 _11803_ (.A(_04295_),
    .B(net3450),
    .Y(_05708_));
 sky130_fd_sc_hd__or2_1 _11804_ (.A(_04506_),
    .B(_04560_),
    .X(_05709_));
 sky130_fd_sc_hd__and2_1 _11805_ (.A(_04561_),
    .B(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__nand2_1 _11806_ (.A(net3451),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _11807_ (.A(_05706_),
    .B(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__and2_1 _11808_ (.A(_05684_),
    .B(_05686_),
    .X(_05713_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(_05687_),
    .B(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__or2_1 _11810_ (.A(_05708_),
    .B(_05710_),
    .X(_05715_));
 sky130_fd_sc_hd__nand2_1 _11811_ (.A(_05711_),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__or2_1 _11812_ (.A(_05714_),
    .B(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__or2_1 _11813_ (.A(_05706_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__a21oi_2 _11814_ (.A1(_05712_),
    .A2(_05718_),
    .B1(_05704_),
    .Y(_05719_));
 sky130_fd_sc_hd__xor2_2 _11815_ (.A(_05673_),
    .B(_05702_),
    .X(_05720_));
 sky130_fd_sc_hd__a21oi_2 _11816_ (.A1(_05719_),
    .A2(_05720_),
    .B1(_05703_),
    .Y(_05721_));
 sky130_fd_sc_hd__xnor2_1 _11817_ (.A(_05637_),
    .B(_05671_),
    .Y(_05722_));
 sky130_fd_sc_hd__or2_1 _11818_ (.A(_05721_),
    .B(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__o21ai_2 _11819_ (.A1(_05721_),
    .A2(_05722_),
    .B1(_05672_),
    .Y(_05724_));
 sky130_fd_sc_hd__o21ba_1 _11820_ (.A1(_05636_),
    .A2(_05724_),
    .B1_N(_05635_),
    .X(_05725_));
 sky130_fd_sc_hd__a21oi_1 _11821_ (.A1(_05596_),
    .A2(_05725_),
    .B1(_05595_),
    .Y(_05726_));
 sky130_fd_sc_hd__a21bo_1 _11822_ (.A1(_04649_),
    .A2(_04650_),
    .B1_N(_04652_),
    .X(_05727_));
 sky130_fd_sc_hd__a21o_1 _11823_ (.A1(_04633_),
    .A2(_04634_),
    .B1(_04607_),
    .X(_05728_));
 sky130_fd_sc_hd__a211o_1 _11824_ (.A1(_04635_),
    .A2(_04636_),
    .B1(_04638_),
    .C1(_05728_),
    .X(_05729_));
 sky130_fd_sc_hd__xnor2_1 _11825_ (.A(_05727_),
    .B(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__a21oi_1 _11826_ (.A1(_04647_),
    .A2(_04648_),
    .B1(_04593_),
    .Y(_05731_));
 sky130_fd_sc_hd__a21bo_1 _11827_ (.A1(_04642_),
    .A2(_04643_),
    .B1_N(_04645_),
    .X(_05732_));
 sky130_fd_sc_hd__a211oi_4 _11828_ (.A1(_04640_),
    .A2(_04641_),
    .B1(_05732_),
    .C1(_04580_),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_2 _11829_ (.A(_05731_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__xnor2_1 _11830_ (.A(_05730_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__or3b_1 _11831_ (.A(_05238_),
    .B(_05496_),
    .C_N(_05225_),
    .X(_05736_));
 sky130_fd_sc_hd__a21o_1 _11832_ (.A1(_04962_),
    .A2(_04977_),
    .B1(_05217_),
    .X(_05737_));
 sky130_fd_sc_hd__or3b_1 _11833_ (.A(_04667_),
    .B(_04674_),
    .C_N(_04938_),
    .X(_05738_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(_05737_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__xnor2_1 _11835_ (.A(_05736_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__xnor2_1 _11836_ (.A(_05735_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nor2_1 _11837_ (.A(_05524_),
    .B(_05526_),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_1 _11838_ (.A(_05505_),
    .B(_05507_),
    .Y(_05743_));
 sky130_fd_sc_hd__o21a_1 _11839_ (.A1(_05220_),
    .A2(_05497_),
    .B1(_05219_),
    .X(_05744_));
 sky130_fd_sc_hd__a21o_1 _11840_ (.A1(_04959_),
    .A2(_04960_),
    .B1(_04941_),
    .X(_05745_));
 sky130_fd_sc_hd__xnor2_2 _11841_ (.A(_05744_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__xnor2_1 _11842_ (.A(_05743_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__xnor2_1 _11843_ (.A(_05742_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__xnor2_1 _11844_ (.A(net3666),
    .B(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__a21oi_1 _11845_ (.A1(_04571_),
    .A2(_05552_),
    .B1(_05550_),
    .Y(_05750_));
 sky130_fd_sc_hd__o31a_1 _11846_ (.A1(_04303_),
    .A2(_04315_),
    .A3(_04573_),
    .B1(_04307_),
    .X(_05751_));
 sky130_fd_sc_hd__and2b_1 _11847_ (.A_N(_04576_),
    .B(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__nand2b_1 _11848_ (.A_N(_04654_),
    .B(_04656_),
    .Y(_05753_));
 sky130_fd_sc_hd__a21o_1 _11849_ (.A1(_04622_),
    .A2(_04623_),
    .B1(net3730),
    .X(_05754_));
 sky130_fd_sc_hd__a211o_1 _11850_ (.A1(_04624_),
    .A2(_04625_),
    .B1(_04628_),
    .C1(net3731),
    .X(_05755_));
 sky130_fd_sc_hd__a21oi_1 _11851_ (.A1(_04578_),
    .A2(_04631_),
    .B1(_04630_),
    .Y(_05756_));
 sky130_fd_sc_hd__xnor2_1 _11852_ (.A(net3732),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__xnor2_1 _11853_ (.A(_05753_),
    .B(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__xnor2_1 _11854_ (.A(_05752_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__xnor2_1 _11855_ (.A(_05750_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__xnor2_1 _11856_ (.A(_05749_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__xnor2_1 _11857_ (.A(_05726_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(net1229),
    .A1(_05762_),
    .S(net250),
    .X(_00381_));
 sky130_fd_sc_hd__nor2_1 _11859_ (.A(_05596_),
    .B(_05725_),
    .Y(_05763_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_05596_),
    .A2(_05725_),
    .B1(net1247),
    .X(_05764_));
 sky130_fd_sc_hd__a2bb2o_1 _11861_ (.A1_N(_05763_),
    .A2_N(_05764_),
    .B1(net1273),
    .B2(net1247),
    .X(_00380_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(_05635_),
    .B(_05636_),
    .Y(_05765_));
 sky130_fd_sc_hd__nand2_1 _11863_ (.A(_05724_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__o21a_1 _11864_ (.A1(_05724_),
    .A2(_05765_),
    .B1(net37),
    .X(_05767_));
 sky130_fd_sc_hd__a22o_1 _11865_ (.A1(net1293),
    .A2(net1247),
    .B1(_05766_),
    .B2(_05767_),
    .X(_00379_));
 sky130_fd_sc_hd__and2_1 _11866_ (.A(net2564),
    .B(net1247),
    .X(_05768_));
 sky130_fd_sc_hd__nand2_1 _11867_ (.A(net3602),
    .B(net3837),
    .Y(_05769_));
 sky130_fd_sc_hd__a31o_1 _11868_ (.A1(net37),
    .A2(_05723_),
    .A3(_05769_),
    .B1(net2566),
    .X(_00378_));
 sky130_fd_sc_hd__nor2_1 _11869_ (.A(_05719_),
    .B(_05720_),
    .Y(_05770_));
 sky130_fd_sc_hd__a21o_1 _11870_ (.A1(_05719_),
    .A2(_05720_),
    .B1(net35),
    .X(_05771_));
 sky130_fd_sc_hd__a2bb2o_1 _11871_ (.A1_N(_05770_),
    .A2_N(_05771_),
    .B1(net1313),
    .B2(net35),
    .X(_00377_));
 sky130_fd_sc_hd__and3_1 _11872_ (.A(_05704_),
    .B(_05712_),
    .C(_05718_),
    .X(_05772_));
 sky130_fd_sc_hd__or2_1 _11873_ (.A(net35),
    .B(_05719_),
    .X(_05773_));
 sky130_fd_sc_hd__a2bb2o_1 _11874_ (.A1_N(_05772_),
    .A2_N(_05773_),
    .B1(net1305),
    .B2(net35),
    .X(_00376_));
 sky130_fd_sc_hd__and2_1 _11875_ (.A(net2546),
    .B(net35),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_1 _11876_ (.A(_05706_),
    .B(_05717_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21bo_1 _11877_ (.A1(_05718_),
    .A2(_05775_),
    .B1_N(_05711_),
    .X(_05776_));
 sky130_fd_sc_hd__a31o_1 _11878_ (.A1(net37),
    .A2(net3452),
    .A3(_05776_),
    .B1(net2548),
    .X(_00375_));
 sky130_fd_sc_hd__and2_1 _11879_ (.A(net2558),
    .B(net35),
    .X(_05777_));
 sky130_fd_sc_hd__nand2_1 _11880_ (.A(_05714_),
    .B(_05716_),
    .Y(_05778_));
 sky130_fd_sc_hd__a31o_1 _11881_ (.A1(net37),
    .A2(_05717_),
    .A3(net3221),
    .B1(net2560),
    .X(_00374_));
 sky130_fd_sc_hd__xnor2_1 _11882_ (.A(_02634_),
    .B(_02660_),
    .Y(_05779_));
 sky130_fd_sc_hd__o21ai_2 _11883_ (.A1(_02905_),
    .A2(_02922_),
    .B1(_02921_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand3_1 _11884_ (.A(_02923_),
    .B(_05779_),
    .C(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21o_1 _11885_ (.A1(_02923_),
    .A2(_05780_),
    .B1(_05779_),
    .X(_05782_));
 sky130_fd_sc_hd__xnor2_1 _11886_ (.A(_02353_),
    .B(_02380_),
    .Y(_05783_));
 sky130_fd_sc_hd__and3_1 _11887_ (.A(_05781_),
    .B(_05782_),
    .C(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__a21oi_1 _11888_ (.A1(_05781_),
    .A2(_05782_),
    .B1(_05783_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _11889_ (.A(_02919_),
    .B(_02920_),
    .Y(_05786_));
 sky130_fd_sc_hd__and2_1 _11890_ (.A(_02921_),
    .B(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__and3_1 _11891_ (.A(_02635_),
    .B(_02643_),
    .C(_02659_),
    .X(_05788_));
 sky130_fd_sc_hd__nor2_1 _11892_ (.A(_02660_),
    .B(_05788_),
    .Y(_05789_));
 sky130_fd_sc_hd__and2_1 _11893_ (.A(_05787_),
    .B(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__nand2_1 _11894_ (.A(_05787_),
    .B(_05789_),
    .Y(_05791_));
 sky130_fd_sc_hd__nor2_1 _11895_ (.A(_05787_),
    .B(_05789_),
    .Y(_05792_));
 sky130_fd_sc_hd__and3_1 _11896_ (.A(_02354_),
    .B(_02362_),
    .C(_02379_),
    .X(_05793_));
 sky130_fd_sc_hd__or2_1 _11897_ (.A(_02380_),
    .B(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__or3_4 _11898_ (.A(_05790_),
    .B(_05792_),
    .C(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__a211oi_2 _11899_ (.A1(_05791_),
    .A2(_05795_),
    .B1(_05784_),
    .C1(_05785_),
    .Y(_05796_));
 sky130_fd_sc_hd__o211a_1 _11900_ (.A1(_05784_),
    .A2(_05785_),
    .B1(_05791_),
    .C1(_05795_),
    .X(_05797_));
 sky130_fd_sc_hd__xor2_2 _11901_ (.A(_01425_),
    .B(_01453_),
    .X(_05798_));
 sky130_fd_sc_hd__xor2_1 _11902_ (.A(_00917_),
    .B(_00944_),
    .X(_05799_));
 sky130_fd_sc_hd__o21ai_1 _11903_ (.A1(_01172_),
    .A2(_01174_),
    .B1(_01202_),
    .Y(_05800_));
 sky130_fd_sc_hd__nand3_1 _11904_ (.A(_01203_),
    .B(_05799_),
    .C(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__a21o_1 _11905_ (.A1(_01203_),
    .A2(_05800_),
    .B1(_05799_),
    .X(_05802_));
 sky130_fd_sc_hd__and3_1 _11906_ (.A(_05798_),
    .B(_05801_),
    .C(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__a21oi_1 _11907_ (.A1(_05801_),
    .A2(_05802_),
    .B1(_05798_),
    .Y(_05804_));
 sky130_fd_sc_hd__or2_1 _11908_ (.A(_05803_),
    .B(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__nor3_1 _11909_ (.A(_05796_),
    .B(_05797_),
    .C(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21a_1 _11910_ (.A1(_05796_),
    .A2(_05797_),
    .B1(_05805_),
    .X(_05807_));
 sky130_fd_sc_hd__o21ai_2 _11911_ (.A1(_05790_),
    .A2(_05792_),
    .B1(_05794_),
    .Y(_05808_));
 sky130_fd_sc_hd__and3_1 _11912_ (.A(_02907_),
    .B(_02914_),
    .C(_02917_),
    .X(_05809_));
 sky130_fd_sc_hd__a211o_1 _11913_ (.A1(_02643_),
    .A2(_02644_),
    .B1(_02651_),
    .C1(_02658_),
    .X(_05810_));
 sky130_fd_sc_hd__nand2_1 _11914_ (.A(_02659_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__nor3_2 _11915_ (.A(_02918_),
    .B(_05809_),
    .C(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21a_1 _11916_ (.A1(_02918_),
    .A2(_05809_),
    .B1(_05811_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_02363_),
    .B(_02378_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand2_1 _11918_ (.A(_02379_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__or3_2 _11919_ (.A(_05812_),
    .B(_05813_),
    .C(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__inv_2 _11920_ (.A(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__o211ai_4 _11921_ (.A1(_05812_),
    .A2(_05817_),
    .B1(_05795_),
    .C1(_05808_),
    .Y(_05818_));
 sky130_fd_sc_hd__a211o_1 _11922_ (.A1(_05795_),
    .A2(_05808_),
    .B1(_05812_),
    .C1(_05817_),
    .X(_05819_));
 sky130_fd_sc_hd__and2_1 _11923_ (.A(_00918_),
    .B(_00943_),
    .X(_05820_));
 sky130_fd_sc_hd__or2_1 _11924_ (.A(_00944_),
    .B(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__nand2_1 _11925_ (.A(_01176_),
    .B(_01200_),
    .Y(_05822_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_01202_),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__nor2_1 _11927_ (.A(_05821_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__and2_1 _11928_ (.A(_05821_),
    .B(_05823_),
    .X(_05825_));
 sky130_fd_sc_hd__and3_1 _11929_ (.A(_01426_),
    .B(_01435_),
    .C(_01452_),
    .X(_05826_));
 sky130_fd_sc_hd__or2_1 _11930_ (.A(_01453_),
    .B(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__or3_2 _11931_ (.A(_05824_),
    .B(_05825_),
    .C(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__o21ai_2 _11932_ (.A1(_05824_),
    .A2(_05825_),
    .B1(_05827_),
    .Y(_05829_));
 sky130_fd_sc_hd__nand4_4 _11933_ (.A(_05818_),
    .B(_05819_),
    .C(_05828_),
    .D(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a211o_1 _11934_ (.A1(_05818_),
    .A2(_05830_),
    .B1(_05806_),
    .C1(_05807_),
    .X(_05831_));
 sky130_fd_sc_hd__o211ai_2 _11935_ (.A1(_05806_),
    .A2(_05807_),
    .B1(_05818_),
    .C1(_05830_),
    .Y(_05832_));
 sky130_fd_sc_hd__or3b_1 _11936_ (.A(_01992_),
    .B(_02000_),
    .C_N(_02001_),
    .X(_05833_));
 sky130_fd_sc_hd__nand2b_2 _11937_ (.A_N(_02002_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__and2b_1 _11938_ (.A_N(_05824_),
    .B(_05828_),
    .X(_05835_));
 sky130_fd_sc_hd__o21bai_1 _11939_ (.A1(_01699_),
    .A2(_01701_),
    .B1_N(_01728_),
    .Y(_05836_));
 sky130_fd_sc_hd__and2_1 _11940_ (.A(_01729_),
    .B(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__nand2b_1 _11941_ (.A_N(_05835_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__xnor2_1 _11942_ (.A(_05835_),
    .B(_05837_),
    .Y(_05839_));
 sky130_fd_sc_hd__inv_2 _11943_ (.A(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__xnor2_1 _11944_ (.A(_05834_),
    .B(_05839_),
    .Y(_05841_));
 sky130_fd_sc_hd__and3_1 _11945_ (.A(_05831_),
    .B(_05832_),
    .C(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__a21bo_1 _11946_ (.A1(_05832_),
    .A2(_05841_),
    .B1_N(_05831_),
    .X(_05843_));
 sky130_fd_sc_hd__a31o_1 _11947_ (.A1(_01203_),
    .A2(_05799_),
    .A3(_05800_),
    .B1(_05803_),
    .X(_05844_));
 sky130_fd_sc_hd__xor2_1 _11948_ (.A(net3726),
    .B(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__xnor2_1 _11949_ (.A(_05843_),
    .B(net3727),
    .Y(_05846_));
 sky130_fd_sc_hd__o211a_1 _11950_ (.A1(_01684_),
    .A2(_01685_),
    .B1(net2777),
    .C1(_01729_),
    .X(_05847_));
 sky130_fd_sc_hd__nor2_1 _11951_ (.A(_01730_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__and2b_1 _11952_ (.A_N(_02615_),
    .B(_02616_),
    .X(_05849_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_05796_),
    .B(_05806_),
    .Y(_05850_));
 sky130_fd_sc_hd__xnor2_1 _11954_ (.A(_01204_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__xnor2_1 _11955_ (.A(_05849_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__xnor2_1 _11956_ (.A(_05848_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__a21oi_1 _11957_ (.A1(_05831_),
    .A2(_05832_),
    .B1(_05841_),
    .Y(_05854_));
 sky130_fd_sc_hd__a22o_1 _11958_ (.A1(_05818_),
    .A2(_05819_),
    .B1(_05828_),
    .B2(_05829_),
    .X(_05855_));
 sky130_fd_sc_hd__o21ai_2 _11959_ (.A1(_05812_),
    .A2(_05813_),
    .B1(_05815_),
    .Y(_05856_));
 sky130_fd_sc_hd__nor2_1 _11960_ (.A(_02655_),
    .B(_02657_),
    .Y(_05857_));
 sky130_fd_sc_hd__nor2_1 _11961_ (.A(_02658_),
    .B(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__xnor2_1 _11962_ (.A(_02915_),
    .B(_02916_),
    .Y(_05859_));
 sky130_fd_sc_hd__and2_2 _11963_ (.A(_05858_),
    .B(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__nor2_1 _11964_ (.A(_05858_),
    .B(_05859_),
    .Y(_05861_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(_02374_),
    .B(_02376_),
    .Y(_05862_));
 sky130_fd_sc_hd__or2_1 _11966_ (.A(_02377_),
    .B(_05862_),
    .X(_05863_));
 sky130_fd_sc_hd__nor3_2 _11967_ (.A(_05860_),
    .B(_05861_),
    .C(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__inv_2 _11968_ (.A(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__o211ai_4 _11969_ (.A1(_05860_),
    .A2(_05864_),
    .B1(_05816_),
    .C1(_05856_),
    .Y(_05866_));
 sky130_fd_sc_hd__inv_2 _11970_ (.A(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__a211o_1 _11971_ (.A1(_05816_),
    .A2(_05856_),
    .B1(_05860_),
    .C1(_05864_),
    .X(_05868_));
 sky130_fd_sc_hd__o211a_1 _11972_ (.A1(_00925_),
    .A2(_00926_),
    .B1(_00934_),
    .C1(_00940_),
    .X(_05869_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(_01184_),
    .B(_01198_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(_01199_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__nor3_1 _11975_ (.A(_00941_),
    .B(_05869_),
    .C(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21a_1 _11976_ (.A1(_00941_),
    .A2(_05869_),
    .B1(_05871_),
    .X(_05873_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(_01436_),
    .B(_01451_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(_01452_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__or3_2 _11979_ (.A(_05872_),
    .B(_05873_),
    .C(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__o21ai_2 _11980_ (.A1(_05872_),
    .A2(_05873_),
    .B1(_05875_),
    .Y(_05877_));
 sky130_fd_sc_hd__and4_2 _11981_ (.A(_05866_),
    .B(_05868_),
    .C(_05876_),
    .D(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__o211ai_4 _11982_ (.A1(_05867_),
    .A2(_05878_),
    .B1(_05830_),
    .C1(_05855_),
    .Y(_05879_));
 sky130_fd_sc_hd__a211o_1 _11983_ (.A1(_05830_),
    .A2(_05855_),
    .B1(_05867_),
    .C1(_05878_),
    .X(_05880_));
 sky130_fd_sc_hd__o2bb2a_1 _11984_ (.A1_N(_01994_),
    .A2_N(_01999_),
    .B1(_01992_),
    .B2(_01993_),
    .X(_05881_));
 sky130_fd_sc_hd__nand2b_1 _11985_ (.A_N(_05872_),
    .B(_05876_),
    .Y(_05882_));
 sky130_fd_sc_hd__and2_1 _11986_ (.A(_01702_),
    .B(_01727_),
    .X(_05883_));
 sky130_fd_sc_hd__nor2_1 _11987_ (.A(_01728_),
    .B(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__xnor2_1 _11988_ (.A(_05882_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__or3_2 _11989_ (.A(_02000_),
    .B(_05881_),
    .C(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__o21ai_2 _11990_ (.A1(_02000_),
    .A2(_05881_),
    .B1(_05885_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand4_4 _11991_ (.A(_05879_),
    .B(_05880_),
    .C(_05886_),
    .D(_05887_),
    .Y(_05888_));
 sky130_fd_sc_hd__a211oi_1 _11992_ (.A1(_05879_),
    .A2(_05888_),
    .B1(_05842_),
    .C1(_05854_),
    .Y(_05889_));
 sky130_fd_sc_hd__o211a_1 _11993_ (.A1(_05842_),
    .A2(_05854_),
    .B1(_05879_),
    .C1(_05888_),
    .X(_05890_));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(_05889_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__a21bo_1 _11995_ (.A1(_05882_),
    .A2(_05884_),
    .B1_N(_05886_),
    .X(_05892_));
 sky130_fd_sc_hd__a21o_1 _11996_ (.A1(_05891_),
    .A2(_05892_),
    .B1(_05889_),
    .X(_05893_));
 sky130_fd_sc_hd__xor2_1 _11997_ (.A(_05891_),
    .B(_05892_),
    .X(_05894_));
 sky130_fd_sc_hd__a22o_1 _11998_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05886_),
    .B2(_05887_),
    .X(_05895_));
 sky130_fd_sc_hd__a22oi_4 _11999_ (.A1(_05866_),
    .A2(_05868_),
    .B1(_05876_),
    .B2(_05877_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_2 _12000_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05863_),
    .Y(_05897_));
 sky130_fd_sc_hd__xnor2_1 _12001_ (.A(_02653_),
    .B(_02654_),
    .Y(_05898_));
 sky130_fd_sc_hd__nor2_1 _12002_ (.A(_02908_),
    .B(_02910_),
    .Y(_05899_));
 sky130_fd_sc_hd__or2_1 _12003_ (.A(_02911_),
    .B(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__nor2_2 _12004_ (.A(_05898_),
    .B(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__nor2_1 _12005_ (.A(_02372_),
    .B(_02373_),
    .Y(_05902_));
 sky130_fd_sc_hd__nor2_1 _12006_ (.A(_02374_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__and2_1 _12007_ (.A(_05898_),
    .B(_05900_),
    .X(_05904_));
 sky130_fd_sc_hd__nor2_1 _12008_ (.A(_05901_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__and2_2 _12009_ (.A(_05903_),
    .B(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__o211ai_4 _12010_ (.A1(_05901_),
    .A2(_05906_),
    .B1(_05865_),
    .C1(_05897_),
    .Y(_05907_));
 sky130_fd_sc_hd__a211o_1 _12011_ (.A1(_05865_),
    .A2(_05897_),
    .B1(_05901_),
    .C1(_05906_),
    .X(_05908_));
 sky130_fd_sc_hd__nor2_1 _12012_ (.A(_01447_),
    .B(_01449_),
    .Y(_05909_));
 sky130_fd_sc_hd__nor2_1 _12013_ (.A(_01450_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__or2_1 _12014_ (.A(_00937_),
    .B(_00939_),
    .X(_05911_));
 sky130_fd_sc_hd__nand2_1 _12015_ (.A(_00940_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__xnor2_1 _12016_ (.A(_01195_),
    .B(_01197_),
    .Y(_05913_));
 sky130_fd_sc_hd__or2_2 _12017_ (.A(_05912_),
    .B(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__nand2_1 _12018_ (.A(_05912_),
    .B(_05913_),
    .Y(_05915_));
 sky130_fd_sc_hd__nand3_2 _12019_ (.A(_05910_),
    .B(_05914_),
    .C(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__a21o_1 _12020_ (.A1(_05914_),
    .A2(_05915_),
    .B1(_05910_),
    .X(_05917_));
 sky130_fd_sc_hd__and4_1 _12021_ (.A(_05907_),
    .B(_05908_),
    .C(_05916_),
    .D(_05917_),
    .X(_05918_));
 sky130_fd_sc_hd__nand4_2 _12022_ (.A(_05907_),
    .B(_05908_),
    .C(_05916_),
    .D(_05917_),
    .Y(_05919_));
 sky130_fd_sc_hd__a211oi_4 _12023_ (.A1(_05907_),
    .A2(_05919_),
    .B1(_05878_),
    .C1(_05896_),
    .Y(_05920_));
 sky130_fd_sc_hd__o211a_1 _12024_ (.A1(_05878_),
    .A2(_05896_),
    .B1(_05907_),
    .C1(_05919_),
    .X(_05921_));
 sky130_fd_sc_hd__xnor2_1 _12025_ (.A(_01994_),
    .B(_01999_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand3_1 _12026_ (.A(_01711_),
    .B(_01718_),
    .C(_01725_),
    .Y(_05923_));
 sky130_fd_sc_hd__nand2_2 _12027_ (.A(_01726_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__a21oi_2 _12028_ (.A1(_05914_),
    .A2(_05916_),
    .B1(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__and3_1 _12029_ (.A(_05914_),
    .B(_05916_),
    .C(_05924_),
    .X(_05926_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(_05925_),
    .B(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__nor2_1 _12031_ (.A(_05922_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__and2_1 _12032_ (.A(_05922_),
    .B(_05927_),
    .X(_05929_));
 sky130_fd_sc_hd__or2_1 _12033_ (.A(_05928_),
    .B(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__nor3_2 _12034_ (.A(_05920_),
    .B(_05921_),
    .C(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__o211ai_2 _12035_ (.A1(_05920_),
    .A2(_05931_),
    .B1(_05888_),
    .C1(_05895_),
    .Y(_05932_));
 sky130_fd_sc_hd__a211o_1 _12036_ (.A1(_05888_),
    .A2(_05895_),
    .B1(_05920_),
    .C1(_05931_),
    .X(_05933_));
 sky130_fd_sc_hd__o211ai_2 _12037_ (.A1(_05925_),
    .A2(_05928_),
    .B1(_05932_),
    .C1(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand2_1 _12038_ (.A(_05932_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand2_1 _12039_ (.A(_05894_),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__xnor2_1 _12040_ (.A(_05894_),
    .B(_05935_),
    .Y(_05937_));
 sky130_fd_sc_hd__a211o_1 _12041_ (.A1(_05932_),
    .A2(_05933_),
    .B1(_05925_),
    .C1(_05928_),
    .X(_05938_));
 sky130_fd_sc_hd__o21a_1 _12042_ (.A1(_05920_),
    .A2(_05921_),
    .B1(_05930_),
    .X(_05939_));
 sky130_fd_sc_hd__a22oi_2 _12043_ (.A1(_05907_),
    .A2(_05908_),
    .B1(_05916_),
    .B2(_05917_),
    .Y(_05940_));
 sky130_fd_sc_hd__nor2_1 _12044_ (.A(_05903_),
    .B(_05905_),
    .Y(_05941_));
 sky130_fd_sc_hd__a22oi_1 _12045_ (.A1(net1648),
    .A2(net2045),
    .B1(net959),
    .B2(net105),
    .Y(_05942_));
 sky130_fd_sc_hd__a22o_1 _12046_ (.A1(net1640),
    .A2(net785),
    .B1(net1725),
    .B2(net1829),
    .X(_05943_));
 sky130_fd_sc_hd__or4b_2 _12047_ (.A(_02654_),
    .B(_02910_),
    .C(_05942_),
    .D_N(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__a2bb2o_1 _12048_ (.A1_N(_02654_),
    .A2_N(_05942_),
    .B1(_05943_),
    .B2(_02909_),
    .X(_05945_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__a22oi_1 _12050_ (.A1(net1603),
    .A2(net2682),
    .B1(net905),
    .B2(net884),
    .Y(_05947_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_02373_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__or3_1 _12052_ (.A(_02373_),
    .B(_05946_),
    .C(_05947_),
    .X(_05949_));
 sky130_fd_sc_hd__a211o_2 _12053_ (.A1(_05944_),
    .A2(_05949_),
    .B1(_05906_),
    .C1(_05941_),
    .X(_05950_));
 sky130_fd_sc_hd__a21oi_1 _12054_ (.A1(_00933_),
    .A2(_00935_),
    .B1(_00936_),
    .Y(_05951_));
 sky130_fd_sc_hd__or2_1 _12055_ (.A(_00937_),
    .B(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__nor2_1 _12056_ (.A(_01193_),
    .B(_01194_),
    .Y(_05953_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(_01195_),
    .B(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__or2_1 _12058_ (.A(_05952_),
    .B(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2_1 _12059_ (.A(_05952_),
    .B(_05954_),
    .Y(_05956_));
 sky130_fd_sc_hd__and2_1 _12060_ (.A(_05955_),
    .B(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__nor2_1 _12061_ (.A(_01445_),
    .B(_01446_),
    .Y(_05958_));
 sky130_fd_sc_hd__nor2_1 _12062_ (.A(_01447_),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2_1 _12063_ (.A(_05957_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(_05957_),
    .B(_05959_),
    .X(_05961_));
 sky130_fd_sc_hd__o211ai_2 _12065_ (.A1(_05906_),
    .A2(_05941_),
    .B1(_05944_),
    .C1(_05949_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand4_2 _12066_ (.A(_05950_),
    .B(_05960_),
    .C(_05961_),
    .D(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a211o_1 _12067_ (.A1(_05950_),
    .A2(_05963_),
    .B1(_05918_),
    .C1(_05940_),
    .X(_05964_));
 sky130_fd_sc_hd__o211ai_2 _12068_ (.A1(_05918_),
    .A2(_05940_),
    .B1(_05950_),
    .C1(_05963_),
    .Y(_05965_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_01995_),
    .B(_01998_),
    .Y(_05966_));
 sky130_fd_sc_hd__or2_1 _12070_ (.A(_01999_),
    .B(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_1 _12071_ (.A(_01722_),
    .B(_01724_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_1 _12072_ (.A(_01725_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__a21o_1 _12073_ (.A1(_05955_),
    .A2(_05960_),
    .B1(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__nand3_1 _12074_ (.A(_05955_),
    .B(_05960_),
    .C(_05969_),
    .Y(_05971_));
 sky130_fd_sc_hd__nand2_1 _12075_ (.A(_05970_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__or2_1 _12076_ (.A(_05967_),
    .B(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__nand2_1 _12077_ (.A(_05967_),
    .B(_05972_),
    .Y(_05974_));
 sky130_fd_sc_hd__and2_1 _12078_ (.A(_05973_),
    .B(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__nand3_2 _12079_ (.A(_05964_),
    .B(_05965_),
    .C(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__a211oi_2 _12080_ (.A1(_05964_),
    .A2(_05976_),
    .B1(_05931_),
    .C1(_05939_),
    .Y(_05977_));
 sky130_fd_sc_hd__o211a_1 _12081_ (.A1(_05931_),
    .A2(_05939_),
    .B1(_05964_),
    .C1(_05976_),
    .X(_05978_));
 sky130_fd_sc_hd__a211oi_2 _12082_ (.A1(_05970_),
    .A2(_05973_),
    .B1(_05977_),
    .C1(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__o211a_1 _12083_ (.A1(_05977_),
    .A2(_05979_),
    .B1(_05934_),
    .C1(_05938_),
    .X(_05980_));
 sky130_fd_sc_hd__a211o_1 _12084_ (.A1(_05934_),
    .A2(_05938_),
    .B1(_05977_),
    .C1(_05979_),
    .X(_05981_));
 sky130_fd_sc_hd__nand2b_1 _12085_ (.A_N(_05980_),
    .B(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__o211a_1 _12086_ (.A1(_05977_),
    .A2(_05978_),
    .B1(_05970_),
    .C1(_05973_),
    .X(_05983_));
 sky130_fd_sc_hd__nor2_1 _12087_ (.A(_05979_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__a21o_1 _12088_ (.A1(_05964_),
    .A2(_05965_),
    .B1(_05975_),
    .X(_05985_));
 sky130_fd_sc_hd__a22o_1 _12089_ (.A1(_05960_),
    .A2(_05961_),
    .B1(_05962_),
    .B2(_05950_),
    .X(_05986_));
 sky130_fd_sc_hd__xnor2_1 _12090_ (.A(_05946_),
    .B(_05948_),
    .Y(_05987_));
 sky130_fd_sc_hd__and4_1 _12091_ (.A(net1640),
    .B(net1648),
    .C(net1725),
    .D(net959),
    .X(_05988_));
 sky130_fd_sc_hd__a22oi_1 _12092_ (.A1(net1640),
    .A2(net1725),
    .B1(net2095),
    .B2(net1648),
    .Y(_05989_));
 sky130_fd_sc_hd__and4bb_1 _12093_ (.A_N(_05988_),
    .B_N(_05989_),
    .C(net1603),
    .D(net905),
    .X(_05990_));
 sky130_fd_sc_hd__nor2_1 _12094_ (.A(_05988_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__and2b_1 _12095_ (.A_N(_05991_),
    .B(_05987_),
    .X(_05992_));
 sky130_fd_sc_hd__xnor2_1 _12096_ (.A(_05987_),
    .B(_05991_),
    .Y(_05993_));
 sky130_fd_sc_hd__inv_2 _12097_ (.A(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__a22oi_1 _12098_ (.A1(net81),
    .A2(net1950),
    .B1(net3724),
    .B2(net887),
    .Y(_05995_));
 sky130_fd_sc_hd__nor2_1 _12099_ (.A(_01446_),
    .B(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__inv_2 _12100_ (.A(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__a22oi_2 _12101_ (.A1(net1644),
    .A2(net764),
    .B1(net2041),
    .B2(net806),
    .Y(_05998_));
 sky130_fd_sc_hd__a22o_1 _12102_ (.A1(net88),
    .A2(net153),
    .B1(net1913),
    .B2(net2136),
    .X(_05999_));
 sky130_fd_sc_hd__inv_2 _12103_ (.A(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__nor4_1 _12104_ (.A(_00936_),
    .B(_01194_),
    .C(_05998_),
    .D(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__o22a_1 _12105_ (.A1(_00936_),
    .A2(_05998_),
    .B1(_06000_),
    .B2(_01194_),
    .X(_06002_));
 sky130_fd_sc_hd__nor2_1 _12106_ (.A(_06001_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__xnor2_1 _12107_ (.A(_05996_),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__nor2_1 _12108_ (.A(_05994_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__o211a_1 _12109_ (.A1(_05992_),
    .A2(_06005_),
    .B1(_05963_),
    .C1(_05986_),
    .X(_06006_));
 sky130_fd_sc_hd__inv_2 _12110_ (.A(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__o21bai_2 _12111_ (.A1(_05997_),
    .A2(_06002_),
    .B1_N(_06001_),
    .Y(_06008_));
 sky130_fd_sc_hd__nor2_1 _12112_ (.A(_01719_),
    .B(_01720_),
    .Y(_06009_));
 sky130_fd_sc_hd__nor2_1 _12113_ (.A(_01721_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__and2_1 _12114_ (.A(_06008_),
    .B(_06010_),
    .X(_06011_));
 sky130_fd_sc_hd__xnor2_1 _12115_ (.A(_06008_),
    .B(_06010_),
    .Y(_06012_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(_01981_),
    .A2(_01996_),
    .B1(_01997_),
    .Y(_06013_));
 sky130_fd_sc_hd__or2_1 _12117_ (.A(_01998_),
    .B(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__nor2_1 _12118_ (.A(_06012_),
    .B(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__and2_1 _12119_ (.A(_06012_),
    .B(_06014_),
    .X(_06016_));
 sky130_fd_sc_hd__a211o_1 _12120_ (.A1(_05963_),
    .A2(_05986_),
    .B1(_05992_),
    .C1(_06005_),
    .X(_06017_));
 sky130_fd_sc_hd__or4b_4 _12121_ (.A(_06006_),
    .B(_06015_),
    .C(_06016_),
    .D_N(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__inv_2 _12122_ (.A(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__o211ai_2 _12123_ (.A1(_06006_),
    .A2(_06019_),
    .B1(_05976_),
    .C1(_05985_),
    .Y(_06020_));
 sky130_fd_sc_hd__a211o_1 _12124_ (.A1(_05976_),
    .A2(_05985_),
    .B1(_06006_),
    .C1(_06019_),
    .X(_06021_));
 sky130_fd_sc_hd__o211ai_2 _12125_ (.A1(_06011_),
    .A2(_06015_),
    .B1(_06020_),
    .C1(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_1 _12126_ (.A(_06020_),
    .B(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__a211o_1 _12127_ (.A1(_06020_),
    .A2(_06021_),
    .B1(_06011_),
    .C1(_06015_),
    .X(_06024_));
 sky130_fd_sc_hd__a2bb2o_1 _12128_ (.A1_N(_06015_),
    .A2_N(_06016_),
    .B1(_06017_),
    .B2(_06007_),
    .X(_06025_));
 sky130_fd_sc_hd__and2_1 _12129_ (.A(_05994_),
    .B(_06004_),
    .X(_06026_));
 sky130_fd_sc_hd__o2bb2a_1 _12130_ (.A1_N(net1603),
    .A2_N(net905),
    .B1(_05988_),
    .B2(_05989_),
    .X(_06027_));
 sky130_fd_sc_hd__nor2_1 _12131_ (.A(_05990_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a22o_1 _12132_ (.A1(net88),
    .A2(net1913),
    .B1(net2041),
    .B2(net1644),
    .X(_06029_));
 sky130_fd_sc_hd__inv_2 _12133_ (.A(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__and4_1 _12134_ (.A(net88),
    .B(net1644),
    .C(net1913),
    .D(net2041),
    .X(_06031_));
 sky130_fd_sc_hd__o2bb2a_1 _12135_ (.A1_N(net81),
    .A2_N(net890),
    .B1(_06030_),
    .B2(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__and4b_1 _12136_ (.A_N(_06031_),
    .B(net890),
    .C(net81),
    .D(_06029_),
    .X(_06033_));
 sky130_fd_sc_hd__nor2_1 _12137_ (.A(_06032_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _12138_ (.A(_06028_),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__nor3_1 _12139_ (.A(_06005_),
    .B(_06026_),
    .C(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__o21a_1 _12140_ (.A1(_06005_),
    .A2(_06026_),
    .B1(_06035_),
    .X(_06037_));
 sky130_fd_sc_hd__or2_1 _12141_ (.A(_06036_),
    .B(_06037_),
    .X(_06038_));
 sky130_fd_sc_hd__a22oi_1 _12142_ (.A1(net1636),
    .A2(net749),
    .B1(net139),
    .B2(net1946),
    .Y(_06039_));
 sky130_fd_sc_hd__or2_1 _12143_ (.A(_01997_),
    .B(_06039_),
    .X(_06040_));
 sky130_fd_sc_hd__a31o_1 _12144_ (.A1(net1309),
    .A2(net890),
    .A3(_06029_),
    .B1(_06031_),
    .X(_06041_));
 sky130_fd_sc_hd__a22oi_1 _12145_ (.A1(net761),
    .A2(net815),
    .B1(net1118),
    .B2(net740),
    .Y(_06042_));
 sky130_fd_sc_hd__nor2_1 _12146_ (.A(_01720_),
    .B(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_06041_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(_06041_),
    .B(_06043_),
    .X(_06045_));
 sky130_fd_sc_hd__nand2_1 _12149_ (.A(_06044_),
    .B(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__or2_1 _12150_ (.A(_06040_),
    .B(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__nand2_1 _12151_ (.A(_06040_),
    .B(_06046_),
    .Y(_06048_));
 sky130_fd_sc_hd__and2_1 _12152_ (.A(_06047_),
    .B(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__and2b_1 _12153_ (.A_N(_06038_),
    .B(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__o211a_1 _12154_ (.A1(_06036_),
    .A2(_06050_),
    .B1(_06018_),
    .C1(_06025_),
    .X(_06051_));
 sky130_fd_sc_hd__a211oi_1 _12155_ (.A1(_06018_),
    .A2(_06025_),
    .B1(_06036_),
    .C1(_06050_),
    .Y(_06052_));
 sky130_fd_sc_hd__or2_1 _12156_ (.A(_06051_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__a21oi_2 _12157_ (.A1(_06044_),
    .A2(_06047_),
    .B1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__o211ai_2 _12158_ (.A1(_06051_),
    .A2(_06054_),
    .B1(_06022_),
    .C1(_06024_),
    .Y(_06055_));
 sky130_fd_sc_hd__and3_1 _12159_ (.A(_06044_),
    .B(_06047_),
    .C(_06053_),
    .X(_06056_));
 sky130_fd_sc_hd__xnor2_1 _12160_ (.A(_06038_),
    .B(_06049_),
    .Y(_06057_));
 sky130_fd_sc_hd__and4_1 _12161_ (.A(net1636),
    .B(net761),
    .C(net139),
    .D(net1118),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__or2_1 _12163_ (.A(_06028_),
    .B(_06034_),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_06035_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__a22oi_2 _12165_ (.A1(net1636),
    .A2(net139),
    .B1(net1118),
    .B2(net761),
    .Y(_06062_));
 sky130_fd_sc_hd__nor3_1 _12166_ (.A(_06058_),
    .B(_06061_),
    .C(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_1 _12167_ (.A(_06057_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__a211oi_4 _12168_ (.A1(net3188),
    .A2(_06064_),
    .B1(_06054_),
    .C1(_06056_),
    .Y(_06065_));
 sky130_fd_sc_hd__a211o_1 _12169_ (.A1(_06022_),
    .A2(_06024_),
    .B1(_06051_),
    .C1(_06054_),
    .X(_06066_));
 sky130_fd_sc_hd__nand3_2 _12170_ (.A(_06055_),
    .B(_06065_),
    .C(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__xnor2_1 _12171_ (.A(_05984_),
    .B(_06023_),
    .Y(_06068_));
 sky130_fd_sc_hd__a21o_1 _12172_ (.A1(_06055_),
    .A2(_06067_),
    .B1(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__a21bo_1 _12173_ (.A1(_05984_),
    .A2(_06023_),
    .B1_N(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__a21oi_2 _12174_ (.A1(_05981_),
    .A2(_06070_),
    .B1(_05980_),
    .Y(_06071_));
 sky130_fd_sc_hd__o21ai_1 _12175_ (.A1(_05937_),
    .A2(_06071_),
    .B1(_05936_),
    .Y(_06072_));
 sky130_fd_sc_hd__xnor2_1 _12176_ (.A(_05893_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__xnor2_2 _12177_ (.A(_02883_),
    .B(_02924_),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_1 _12178_ (.A(_01154_),
    .B(_01156_),
    .Y(_06075_));
 sky130_fd_sc_hd__o21a_1 _12179_ (.A1(_05834_),
    .A2(_05840_),
    .B1(_05838_),
    .X(_06076_));
 sky130_fd_sc_hd__xnor2_1 _12180_ (.A(_02661_),
    .B(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__xnor2_2 _12181_ (.A(_01407_),
    .B(_01454_),
    .Y(_06078_));
 sky130_fd_sc_hd__nor2_1 _12182_ (.A(_00896_),
    .B(_00897_),
    .Y(_06079_));
 sky130_fd_sc_hd__and2b_1 _12183_ (.A_N(_02334_),
    .B(_02335_),
    .X(_06080_));
 sky130_fd_sc_hd__xnor2_1 _12184_ (.A(_06079_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__xnor2_1 _12185_ (.A(_06078_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__xnor2_1 _12186_ (.A(_06077_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__xor2_1 _12187_ (.A(_06075_),
    .B(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__xnor2_1 _12188_ (.A(_06074_),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__xnor2_1 _12189_ (.A(_06073_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__xnor2_1 _12190_ (.A(net3745),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nor3_1 _12191_ (.A(_01951_),
    .B(_01973_),
    .C(_02002_),
    .Y(_06088_));
 sky130_fd_sc_hd__nor2_1 _12192_ (.A(_02003_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a31o_1 _12193_ (.A1(_02923_),
    .A2(_05779_),
    .A3(_05780_),
    .B1(_05784_),
    .X(_06090_));
 sky130_fd_sc_hd__xor2_1 _12194_ (.A(_02381_),
    .B(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__xor2_1 _12195_ (.A(_06089_),
    .B(net3672),
    .X(_06092_));
 sky130_fd_sc_hd__xnor2_1 _12196_ (.A(_06087_),
    .B(net3673),
    .Y(_06093_));
 sky130_fd_sc_hd__xnor2_1 _12197_ (.A(net3728),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(net1289),
    .A1(_06094_),
    .S(net37),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(_05937_),
    .B(_06071_),
    .Y(_06095_));
 sky130_fd_sc_hd__o21a_1 _12200_ (.A1(_05937_),
    .A2(_06071_),
    .B1(net37),
    .X(_06096_));
 sky130_fd_sc_hd__a22o_1 _12201_ (.A1(net1285),
    .A2(net34),
    .B1(_06095_),
    .B2(_06096_),
    .X(_00372_));
 sky130_fd_sc_hd__xnor2_1 _12202_ (.A(_05982_),
    .B(_06070_),
    .Y(_06097_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(net1269),
    .A1(_06097_),
    .S(net37),
    .X(_00371_));
 sky130_fd_sc_hd__and3_1 _12204_ (.A(_06055_),
    .B(_06067_),
    .C(_06068_),
    .X(_06098_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(net37),
    .B(_06069_),
    .Y(_06099_));
 sky130_fd_sc_hd__a2bb2o_1 _12206_ (.A1_N(_06098_),
    .A2_N(_06099_),
    .B1(net1251),
    .B2(net34),
    .X(_00370_));
 sky130_fd_sc_hd__and2_1 _12207_ (.A(net1415),
    .B(net34),
    .X(_06100_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(_06055_),
    .A2(_06066_),
    .B1(_06065_),
    .X(_06101_));
 sky130_fd_sc_hd__a31o_1 _12209_ (.A1(net37),
    .A2(net3190),
    .A3(_06101_),
    .B1(net1417),
    .X(_00369_));
 sky130_fd_sc_hd__o211a_1 _12210_ (.A1(_06054_),
    .A2(_06056_),
    .B1(_06059_),
    .C1(_06064_),
    .X(_06102_));
 sky130_fd_sc_hd__or3_1 _12211_ (.A(net34),
    .B(_06065_),
    .C(_06102_),
    .X(_06103_));
 sky130_fd_sc_hd__a21bo_1 _12212_ (.A1(net1211),
    .A2(net1247),
    .B1_N(_06103_),
    .X(_00368_));
 sky130_fd_sc_hd__or2_1 _12213_ (.A(_06057_),
    .B(_06063_),
    .X(_06104_));
 sky130_fd_sc_hd__and2_1 _12214_ (.A(_06064_),
    .B(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__o211a_1 _12215_ (.A1(_06058_),
    .A2(_06105_),
    .B1(_06059_),
    .C1(net37),
    .X(_06106_));
 sky130_fd_sc_hd__a21o_1 _12216_ (.A1(net1225),
    .A2(net36),
    .B1(_06106_),
    .X(_00367_));
 sky130_fd_sc_hd__o21a_1 _12217_ (.A1(_06058_),
    .A2(_06062_),
    .B1(_06061_),
    .X(_06107_));
 sky130_fd_sc_hd__or2_1 _12218_ (.A(net34),
    .B(_06063_),
    .X(_06108_));
 sky130_fd_sc_hd__a2bb2o_1 _12219_ (.A1_N(_06107_),
    .A2_N(_06108_),
    .B1(net1188),
    .B2(net34),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_2 _12220_ (.A(_03491_),
    .B(_03517_),
    .Y(_06109_));
 sky130_fd_sc_hd__xnor2_1 _12221_ (.A(_03744_),
    .B(_03770_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand2_1 _12222_ (.A(_06109_),
    .B(_06110_),
    .Y(_06111_));
 sky130_fd_sc_hd__xor2_2 _12223_ (.A(_03996_),
    .B(_04022_),
    .X(_06112_));
 sky130_fd_sc_hd__or2_1 _12224_ (.A(_06109_),
    .B(_06110_),
    .X(_06113_));
 sky130_fd_sc_hd__and3_1 _12225_ (.A(_06111_),
    .B(_06112_),
    .C(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__a21o_1 _12226_ (.A1(_06109_),
    .A2(_06110_),
    .B1(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__a21oi_1 _12227_ (.A1(_04913_),
    .A2(_04926_),
    .B1(_04925_),
    .Y(_06116_));
 sky130_fd_sc_hd__or2_1 _12228_ (.A(_04927_),
    .B(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__xnor2_2 _12229_ (.A(_05180_),
    .B(_05207_),
    .Y(_06118_));
 sky130_fd_sc_hd__xnor2_1 _12230_ (.A(_06117_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__xor2_2 _12231_ (.A(_05462_),
    .B(_05486_),
    .X(_06120_));
 sky130_fd_sc_hd__nand2b_1 _12232_ (.A_N(_06119_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__xnor2_1 _12233_ (.A(_06119_),
    .B(_06120_),
    .Y(_06122_));
 sky130_fd_sc_hd__a21oi_1 _12234_ (.A1(_04912_),
    .A2(_04924_),
    .B1(_04923_),
    .Y(_06123_));
 sky130_fd_sc_hd__or2_1 _12235_ (.A(_04925_),
    .B(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__and3_1 _12236_ (.A(_05181_),
    .B(_05189_),
    .C(_05206_),
    .X(_06125_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(_05207_),
    .B(_06125_),
    .X(_06126_));
 sky130_fd_sc_hd__nor2_1 _12238_ (.A(_06124_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__and2_1 _12239_ (.A(_06124_),
    .B(_06126_),
    .X(_06128_));
 sky130_fd_sc_hd__or2_1 _12240_ (.A(_06127_),
    .B(_06128_),
    .X(_06129_));
 sky130_fd_sc_hd__nor2_1 _12241_ (.A(_05470_),
    .B(_05471_),
    .Y(_06130_));
 sky130_fd_sc_hd__xnor2_1 _12242_ (.A(_05485_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__o21ba_1 _12243_ (.A1(_06129_),
    .A2(_06131_),
    .B1_N(_06127_),
    .X(_06132_));
 sky130_fd_sc_hd__and2b_1 _12244_ (.A_N(_06132_),
    .B(_06122_),
    .X(_06133_));
 sky130_fd_sc_hd__xnor2_1 _12245_ (.A(_06122_),
    .B(_06132_),
    .Y(_06134_));
 sky130_fd_sc_hd__a21oi_1 _12246_ (.A1(_06111_),
    .A2(_06113_),
    .B1(_06112_),
    .Y(_06135_));
 sky130_fd_sc_hd__nor2_1 _12247_ (.A(_06114_),
    .B(_06135_),
    .Y(_06136_));
 sky130_fd_sc_hd__xnor2_1 _12248_ (.A(_06134_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__xnor2_1 _12249_ (.A(_06129_),
    .B(_06131_),
    .Y(_06138_));
 sky130_fd_sc_hd__nor2_1 _12250_ (.A(_04914_),
    .B(_04922_),
    .Y(_06139_));
 sky130_fd_sc_hd__or2_1 _12251_ (.A(_04923_),
    .B(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__nand2_1 _12252_ (.A(_05190_),
    .B(_05205_),
    .Y(_06141_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_05206_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__or2_1 _12254_ (.A(_06140_),
    .B(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(_06140_),
    .B(_06142_),
    .Y(_06144_));
 sky130_fd_sc_hd__xnor2_1 _12256_ (.A(_05479_),
    .B(_05483_),
    .Y(_06145_));
 sky130_fd_sc_hd__and3_1 _12257_ (.A(_06143_),
    .B(_06144_),
    .C(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__inv_2 _12258_ (.A(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__a21o_1 _12259_ (.A1(_06143_),
    .A2(_06147_),
    .B1(_06138_),
    .X(_06148_));
 sky130_fd_sc_hd__nand3_1 _12260_ (.A(_06138_),
    .B(_06143_),
    .C(_06147_),
    .Y(_06149_));
 sky130_fd_sc_hd__and2_1 _12261_ (.A(_03492_),
    .B(_03516_),
    .X(_06150_));
 sky130_fd_sc_hd__nor2_1 _12262_ (.A(_03517_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__and3_1 _12263_ (.A(_03745_),
    .B(_03753_),
    .C(_03769_),
    .X(_06152_));
 sky130_fd_sc_hd__nor2_1 _12264_ (.A(_03770_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__and2_1 _12265_ (.A(_06151_),
    .B(_06153_),
    .X(_06154_));
 sky130_fd_sc_hd__nor2_1 _12266_ (.A(_06151_),
    .B(_06153_),
    .Y(_06155_));
 sky130_fd_sc_hd__nor2_1 _12267_ (.A(_06154_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__and3_1 _12268_ (.A(_03997_),
    .B(_04004_),
    .C(_04021_),
    .X(_06157_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(_04022_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__and2_1 _12270_ (.A(_06156_),
    .B(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__nor2_1 _12271_ (.A(_06156_),
    .B(_06158_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_1 _12272_ (.A(_06159_),
    .B(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__nand3_2 _12273_ (.A(_06148_),
    .B(_06149_),
    .C(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__a21oi_1 _12274_ (.A1(_06148_),
    .A2(_06162_),
    .B1(_06137_),
    .Y(_06163_));
 sky130_fd_sc_hd__and3_1 _12275_ (.A(_06137_),
    .B(_06148_),
    .C(_06162_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(_06163_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__o21ai_1 _12277_ (.A1(_04264_),
    .A2(_04266_),
    .B1(_04292_),
    .Y(_06166_));
 sky130_fd_sc_hd__and2_1 _12278_ (.A(_04293_),
    .B(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__o21a_1 _12279_ (.A1(_06154_),
    .A2(_06159_),
    .B1(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__nor3_1 _12280_ (.A(_06154_),
    .B(_06159_),
    .C(_06167_),
    .Y(_06169_));
 sky130_fd_sc_hd__or2_1 _12281_ (.A(_06168_),
    .B(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__inv_2 _12282_ (.A(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__or3_1 _12283_ (.A(_04528_),
    .B(_04544_),
    .C(_04558_),
    .X(_06172_));
 sky130_fd_sc_hd__and2_2 _12284_ (.A(_04559_),
    .B(_06172_),
    .X(_06173_));
 sky130_fd_sc_hd__xor2_1 _12285_ (.A(_06170_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__xnor2_1 _12286_ (.A(_06165_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__a21o_1 _12287_ (.A1(_06148_),
    .A2(_06149_),
    .B1(_06161_),
    .X(_06176_));
 sky130_fd_sc_hd__a21oi_1 _12288_ (.A1(_06143_),
    .A2(_06144_),
    .B1(_06145_),
    .Y(_06177_));
 sky130_fd_sc_hd__and2b_1 _12289_ (.A_N(_04921_),
    .B(_04915_),
    .X(_06178_));
 sky130_fd_sc_hd__or2_1 _12290_ (.A(_04922_),
    .B(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__xnor2_1 _12291_ (.A(_05202_),
    .B(_05204_),
    .Y(_06180_));
 sky130_fd_sc_hd__or2_2 _12292_ (.A(_06179_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_06179_),
    .B(_06180_),
    .Y(_06182_));
 sky130_fd_sc_hd__a21bo_1 _12294_ (.A1(_05475_),
    .A2(_05477_),
    .B1_N(_05474_),
    .X(_06183_));
 sky130_fd_sc_hd__xnor2_2 _12295_ (.A(_05472_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand3_4 _12296_ (.A(_06181_),
    .B(_06182_),
    .C(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__a211oi_2 _12297_ (.A1(_06181_),
    .A2(_06185_),
    .B1(_06146_),
    .C1(_06177_),
    .Y(_06186_));
 sky130_fd_sc_hd__o211a_1 _12298_ (.A1(_06146_),
    .A2(_06177_),
    .B1(_06181_),
    .C1(_06185_),
    .X(_06187_));
 sky130_fd_sc_hd__or2_1 _12299_ (.A(_06186_),
    .B(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__xnor2_1 _12300_ (.A(_03501_),
    .B(_03515_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _12301_ (.A(_03754_),
    .B(_03768_),
    .Y(_06190_));
 sky130_fd_sc_hd__nand2_1 _12302_ (.A(_03769_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__or2_1 _12303_ (.A(_06189_),
    .B(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__nand2_1 _12304_ (.A(_06189_),
    .B(_06191_),
    .Y(_06193_));
 sky130_fd_sc_hd__and2_1 _12305_ (.A(_06192_),
    .B(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__inv_2 _12306_ (.A(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__xnor2_2 _12307_ (.A(_04006_),
    .B(_04020_),
    .Y(_06196_));
 sky130_fd_sc_hd__xor2_1 _12308_ (.A(_06194_),
    .B(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(_06188_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__o211ai_2 _12310_ (.A1(_06186_),
    .A2(_06198_),
    .B1(_06162_),
    .C1(_06176_),
    .Y(_06199_));
 sky130_fd_sc_hd__a211o_1 _12311_ (.A1(_06162_),
    .A2(_06176_),
    .B1(_06186_),
    .C1(_06198_),
    .X(_06200_));
 sky130_fd_sc_hd__xnor2_2 _12312_ (.A(_04545_),
    .B(_04557_),
    .Y(_06201_));
 sky130_fd_sc_hd__o21ai_1 _12313_ (.A1(_06195_),
    .A2(_06196_),
    .B1(_06192_),
    .Y(_06202_));
 sky130_fd_sc_hd__nand3_1 _12314_ (.A(_04267_),
    .B(_04274_),
    .C(_04291_),
    .Y(_06203_));
 sky130_fd_sc_hd__and2_1 _12315_ (.A(_04292_),
    .B(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__xor2_1 _12316_ (.A(_06202_),
    .B(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__nand2_1 _12317_ (.A(_06201_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__or2_1 _12318_ (.A(_06201_),
    .B(_06205_),
    .X(_06207_));
 sky130_fd_sc_hd__and2_1 _12319_ (.A(_06206_),
    .B(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__nand3_1 _12320_ (.A(_06199_),
    .B(_06200_),
    .C(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__nand2_1 _12321_ (.A(_06199_),
    .B(_06209_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _12322_ (.A(_06175_),
    .B(_06210_),
    .Y(_06211_));
 sky130_fd_sc_hd__a21bo_1 _12323_ (.A1(_06202_),
    .A2(_06204_),
    .B1_N(_06206_),
    .X(_06212_));
 sky130_fd_sc_hd__and2b_1 _12324_ (.A_N(_06211_),
    .B(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a21oi_1 _12325_ (.A1(_06175_),
    .A2(_06210_),
    .B1(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__xnor2_1 _12326_ (.A(_06115_),
    .B(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__a21oi_1 _12327_ (.A1(_06171_),
    .A2(_06173_),
    .B1(_06168_),
    .Y(_06216_));
 sky130_fd_sc_hd__xnor2_1 _12328_ (.A(_05208_),
    .B(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__xnor2_1 _12329_ (.A(_03978_),
    .B(_04023_),
    .Y(_06218_));
 sky130_fd_sc_hd__and2b_1 _12330_ (.A_N(_03472_),
    .B(_03473_),
    .X(_06219_));
 sky130_fd_sc_hd__nand2_1 _12331_ (.A(_05426_),
    .B(_05444_),
    .Y(_06220_));
 sky130_fd_sc_hd__and2_1 _12332_ (.A(_05460_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__xnor2_1 _12333_ (.A(_06219_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__xnor2_1 _12334_ (.A(_06218_),
    .B(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__xnor2_1 _12335_ (.A(_06217_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__xnor2_1 _12336_ (.A(_03771_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__xor2_1 _12337_ (.A(_06215_),
    .B(net3677),
    .X(_06226_));
 sky130_fd_sc_hd__o211ai_1 _12338_ (.A1(_04246_),
    .A2(_04248_),
    .B1(_04265_),
    .C1(_04293_),
    .Y(_06227_));
 sky130_fd_sc_hd__nand2_1 _12339_ (.A(_04294_),
    .B(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__and3_1 _12340_ (.A(_04507_),
    .B(_04527_),
    .C(_04559_),
    .X(_06229_));
 sky130_fd_sc_hd__nor2_1 _12341_ (.A(_04560_),
    .B(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__xnor2_1 _12342_ (.A(_06211_),
    .B(_06212_),
    .Y(_06231_));
 sky130_fd_sc_hd__a21o_1 _12343_ (.A1(_06199_),
    .A2(_06200_),
    .B1(_06208_),
    .X(_06232_));
 sky130_fd_sc_hd__xnor2_1 _12344_ (.A(_06188_),
    .B(_06197_),
    .Y(_06233_));
 sky130_fd_sc_hd__a21o_1 _12345_ (.A1(_06181_),
    .A2(_06182_),
    .B1(_06184_),
    .X(_06234_));
 sky130_fd_sc_hd__xor2_1 _12346_ (.A(_04917_),
    .B(_04920_),
    .X(_06235_));
 sky130_fd_sc_hd__inv_2 _12347_ (.A(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__xnor2_1 _12348_ (.A(_05199_),
    .B(_05200_),
    .Y(_06237_));
 sky130_fd_sc_hd__nor2_2 _12349_ (.A(_06236_),
    .B(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__xor2_2 _12350_ (.A(_05476_),
    .B(_05477_),
    .X(_06239_));
 sky130_fd_sc_hd__and2_1 _12351_ (.A(_06236_),
    .B(_06237_),
    .X(_06240_));
 sky130_fd_sc_hd__or2_1 _12352_ (.A(_06238_),
    .B(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__nor2_2 _12353_ (.A(_06239_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__o211ai_4 _12354_ (.A1(_06238_),
    .A2(_06242_),
    .B1(_06185_),
    .C1(_06234_),
    .Y(_06243_));
 sky130_fd_sc_hd__a211o_1 _12355_ (.A1(_06185_),
    .A2(_06234_),
    .B1(_06238_),
    .C1(_06242_),
    .X(_06244_));
 sky130_fd_sc_hd__xor2_2 _12356_ (.A(_04017_),
    .B(_04019_),
    .X(_06245_));
 sky130_fd_sc_hd__xnor2_1 _12357_ (.A(_03512_),
    .B(_03514_),
    .Y(_06246_));
 sky130_fd_sc_hd__xnor2_1 _12358_ (.A(_03765_),
    .B(_03767_),
    .Y(_06247_));
 sky130_fd_sc_hd__or2_1 _12359_ (.A(_06246_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__nand2_1 _12360_ (.A(_06246_),
    .B(_06247_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand3_2 _12361_ (.A(_06245_),
    .B(_06248_),
    .C(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__a21o_1 _12362_ (.A1(_06248_),
    .A2(_06249_),
    .B1(_06245_),
    .X(_06251_));
 sky130_fd_sc_hd__nand4_2 _12363_ (.A(_06243_),
    .B(_06244_),
    .C(_06250_),
    .D(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__a21oi_2 _12364_ (.A1(_06243_),
    .A2(_06252_),
    .B1(_06233_),
    .Y(_06253_));
 sky130_fd_sc_hd__and3_1 _12365_ (.A(_06233_),
    .B(_06243_),
    .C(_06252_),
    .X(_06254_));
 sky130_fd_sc_hd__xnor2_2 _12366_ (.A(_04547_),
    .B(_04556_),
    .Y(_06255_));
 sky130_fd_sc_hd__xnor2_2 _12367_ (.A(_04276_),
    .B(_04290_),
    .Y(_06256_));
 sky130_fd_sc_hd__a21oi_1 _12368_ (.A1(_06248_),
    .A2(_06250_),
    .B1(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__and3_1 _12369_ (.A(_06248_),
    .B(_06250_),
    .C(_06256_),
    .X(_06258_));
 sky130_fd_sc_hd__nor2_1 _12370_ (.A(_06257_),
    .B(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__xnor2_1 _12371_ (.A(_06255_),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__or3_2 _12372_ (.A(_06253_),
    .B(_06254_),
    .C(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__inv_2 _12373_ (.A(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__o211a_1 _12374_ (.A1(_06253_),
    .A2(_06262_),
    .B1(_06209_),
    .C1(_06232_),
    .X(_06263_));
 sky130_fd_sc_hd__a211oi_1 _12375_ (.A1(_06209_),
    .A2(_06232_),
    .B1(_06253_),
    .C1(_06262_),
    .Y(_06264_));
 sky130_fd_sc_hd__or2_1 _12376_ (.A(_06263_),
    .B(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__a21o_1 _12377_ (.A1(_06255_),
    .A2(_06259_),
    .B1(_06257_),
    .X(_06266_));
 sky130_fd_sc_hd__and2b_1 _12378_ (.A_N(_06265_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__o21a_1 _12379_ (.A1(_06263_),
    .A2(_06267_),
    .B1(_06231_),
    .X(_06268_));
 sky130_fd_sc_hd__nor3_1 _12380_ (.A(_06231_),
    .B(_06263_),
    .C(_06267_),
    .Y(_06269_));
 sky130_fd_sc_hd__nor2_1 _12381_ (.A(_06268_),
    .B(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__xnor2_1 _12382_ (.A(_06265_),
    .B(_06266_),
    .Y(_06271_));
 sky130_fd_sc_hd__o21ai_1 _12383_ (.A1(_06253_),
    .A2(_06254_),
    .B1(_06260_),
    .Y(_06272_));
 sky130_fd_sc_hd__a22o_1 _12384_ (.A1(_06243_),
    .A2(_06244_),
    .B1(_06250_),
    .B2(_06251_),
    .X(_06273_));
 sky130_fd_sc_hd__nand2_1 _12385_ (.A(_06252_),
    .B(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__and2_1 _12386_ (.A(_06239_),
    .B(_06241_),
    .X(_06275_));
 sky130_fd_sc_hd__nor2_1 _12387_ (.A(_06242_),
    .B(_06275_),
    .Y(_06276_));
 sky130_fd_sc_hd__a22oi_1 _12388_ (.A1(net1615),
    .A2(net1007),
    .B1(net1010),
    .B2(net1934),
    .Y(_06277_));
 sky130_fd_sc_hd__a22o_1 _12389_ (.A1(net1626),
    .A2(net1954),
    .B1(net2333),
    .B2(net968),
    .X(_06278_));
 sky130_fd_sc_hd__or4b_1 _12390_ (.A(_04916_),
    .B(_05200_),
    .C(_06277_),
    .D_N(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a2bb2o_1 _12391_ (.A1_N(_04916_),
    .A2_N(_06277_),
    .B1(_06278_),
    .B2(_05201_),
    .X(_06280_));
 sky130_fd_sc_hd__nand2_1 _12392_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__a22oi_1 _12393_ (.A1(net1611),
    .A2(net2132),
    .B1(net2239),
    .B2(net1721),
    .Y(_06282_));
 sky130_fd_sc_hd__or2_2 _12394_ (.A(_05477_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__o21ai_2 _12395_ (.A1(_06281_),
    .A2(_06283_),
    .B1(_06279_),
    .Y(_06284_));
 sky130_fd_sc_hd__nand2_2 _12396_ (.A(_06276_),
    .B(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__xnor2_1 _12397_ (.A(_03510_),
    .B(_03511_),
    .Y(_06286_));
 sky130_fd_sc_hd__xnor2_1 _12398_ (.A(_03763_),
    .B(_03764_),
    .Y(_06287_));
 sky130_fd_sc_hd__or2_1 _12399_ (.A(_06286_),
    .B(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__nand2_1 _12400_ (.A(_06286_),
    .B(_06287_),
    .Y(_06289_));
 sky130_fd_sc_hd__and2_1 _12401_ (.A(_06288_),
    .B(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__nor2_1 _12402_ (.A(_04015_),
    .B(_04016_),
    .Y(_06291_));
 sky130_fd_sc_hd__nor2_1 _12403_ (.A(_04017_),
    .B(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_2 _12404_ (.A(_06290_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__or2_1 _12405_ (.A(_06290_),
    .B(_06292_),
    .X(_06294_));
 sky130_fd_sc_hd__or2_1 _12406_ (.A(_06276_),
    .B(_06284_),
    .X(_06295_));
 sky130_fd_sc_hd__nand4_4 _12407_ (.A(_06285_),
    .B(_06293_),
    .C(_06294_),
    .D(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__a21oi_2 _12408_ (.A1(_06285_),
    .A2(_06296_),
    .B1(_06274_),
    .Y(_06297_));
 sky130_fd_sc_hd__and3_1 _12409_ (.A(_06274_),
    .B(_06285_),
    .C(_06296_),
    .X(_06298_));
 sky130_fd_sc_hd__nor2_1 _12410_ (.A(_04548_),
    .B(_04555_),
    .Y(_06299_));
 sky130_fd_sc_hd__nor2_2 _12411_ (.A(_04556_),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__xnor2_2 _12412_ (.A(_04287_),
    .B(_04289_),
    .Y(_06301_));
 sky130_fd_sc_hd__a21oi_1 _12413_ (.A1(_06288_),
    .A2(_06293_),
    .B1(_06301_),
    .Y(_06302_));
 sky130_fd_sc_hd__and3_1 _12414_ (.A(_06288_),
    .B(_06293_),
    .C(_06301_),
    .X(_06303_));
 sky130_fd_sc_hd__nor2_1 _12415_ (.A(_06302_),
    .B(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__xnor2_1 _12416_ (.A(_06300_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__nor3_2 _12417_ (.A(_06297_),
    .B(_06298_),
    .C(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__o211a_1 _12418_ (.A1(_06297_),
    .A2(_06306_),
    .B1(_06261_),
    .C1(_06272_),
    .X(_06307_));
 sky130_fd_sc_hd__a211o_1 _12419_ (.A1(_06261_),
    .A2(_06272_),
    .B1(_06297_),
    .C1(_06306_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2b_1 _12420_ (.A_N(_06307_),
    .B(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__a21o_1 _12421_ (.A1(_06300_),
    .A2(_06304_),
    .B1(_06302_),
    .X(_06310_));
 sky130_fd_sc_hd__a21o_1 _12422_ (.A1(_06308_),
    .A2(_06310_),
    .B1(_06307_),
    .X(_06311_));
 sky130_fd_sc_hd__and2_1 _12423_ (.A(_06271_),
    .B(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__xor2_1 _12424_ (.A(_06271_),
    .B(_06311_),
    .X(_06313_));
 sky130_fd_sc_hd__xnor2_1 _12425_ (.A(_06309_),
    .B(_06310_),
    .Y(_06314_));
 sky130_fd_sc_hd__o21a_1 _12426_ (.A1(_06297_),
    .A2(_06298_),
    .B1(_06305_),
    .X(_06315_));
 sky130_fd_sc_hd__a22o_1 _12427_ (.A1(_06293_),
    .A2(_06294_),
    .B1(_06295_),
    .B2(_06285_),
    .X(_06316_));
 sky130_fd_sc_hd__xor2_2 _12428_ (.A(_06281_),
    .B(_06283_),
    .X(_06317_));
 sky130_fd_sc_hd__and4_1 _12429_ (.A(net1626),
    .B(net1615),
    .C(net2333),
    .D(net1010),
    .X(_06318_));
 sky130_fd_sc_hd__a22oi_1 _12430_ (.A1(net1626),
    .A2(net2333),
    .B1(net1010),
    .B2(net1615),
    .Y(_06319_));
 sky130_fd_sc_hd__and4bb_1 _12431_ (.A_N(_06318_),
    .B_N(_06319_),
    .C(net1611),
    .D(net2239),
    .X(_06320_));
 sky130_fd_sc_hd__nor2_1 _12432_ (.A(_06318_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__and2b_2 _12433_ (.A_N(_06321_),
    .B(_06317_),
    .X(_06322_));
 sky130_fd_sc_hd__xnor2_2 _12434_ (.A(_06317_),
    .B(_06321_),
    .Y(_06323_));
 sky130_fd_sc_hd__inv_2 _12435_ (.A(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__a22oi_1 _12436_ (.A1(net1632),
    .A2(net1767),
    .B1(net821),
    .B2(net1773),
    .Y(_06325_));
 sky130_fd_sc_hd__nor2_1 _12437_ (.A(_04016_),
    .B(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__inv_2 _12438_ (.A(_06326_),
    .Y(_06327_));
 sky130_fd_sc_hd__a22oi_2 _12439_ (.A1(net1590),
    .A2(net1809),
    .B1(net2379),
    .B2(net1677),
    .Y(_06328_));
 sky130_fd_sc_hd__a22o_1 _12440_ (.A1(net1607),
    .A2(net1805),
    .B1(net2078),
    .B2(net1752),
    .X(_06329_));
 sky130_fd_sc_hd__inv_2 _12441_ (.A(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__nor4_1 _12442_ (.A(_03511_),
    .B(_03764_),
    .C(_06328_),
    .D(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__o22a_1 _12443_ (.A1(_03511_),
    .A2(_06328_),
    .B1(_06330_),
    .B2(_03764_),
    .X(_06332_));
 sky130_fd_sc_hd__or2_1 _12444_ (.A(_06331_),
    .B(_06332_),
    .X(_06333_));
 sky130_fd_sc_hd__nor2_1 _12445_ (.A(_06327_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__and2_1 _12446_ (.A(_06327_),
    .B(_06333_),
    .X(_06335_));
 sky130_fd_sc_hd__or2_1 _12447_ (.A(_06334_),
    .B(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nor2_2 _12448_ (.A(_06324_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__o211ai_4 _12449_ (.A1(_06322_),
    .A2(_06337_),
    .B1(_06296_),
    .C1(_06316_),
    .Y(_06338_));
 sky130_fd_sc_hd__inv_2 _12450_ (.A(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor2_1 _12451_ (.A(_04285_),
    .B(_04286_),
    .Y(_06340_));
 sky130_fd_sc_hd__nor2_1 _12452_ (.A(_04287_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__o21a_1 _12453_ (.A1(_06331_),
    .A2(_06334_),
    .B1(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nor3_1 _12454_ (.A(_06331_),
    .B(_06334_),
    .C(_06341_),
    .Y(_06343_));
 sky130_fd_sc_hd__nor2_1 _12455_ (.A(_06342_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__xor2_2 _12456_ (.A(_04551_),
    .B(_04554_),
    .X(_06345_));
 sky130_fd_sc_hd__and2_1 _12457_ (.A(_06344_),
    .B(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__nor2_1 _12458_ (.A(_06344_),
    .B(_06345_),
    .Y(_06347_));
 sky130_fd_sc_hd__a211o_1 _12459_ (.A1(_06296_),
    .A2(_06316_),
    .B1(_06322_),
    .C1(_06337_),
    .X(_06348_));
 sky130_fd_sc_hd__or4b_2 _12460_ (.A(_06339_),
    .B(_06346_),
    .C(_06347_),
    .D_N(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a211o_1 _12461_ (.A1(_06338_),
    .A2(_06349_),
    .B1(_06306_),
    .C1(_06315_),
    .X(_06350_));
 sky130_fd_sc_hd__o211ai_2 _12462_ (.A1(_06306_),
    .A2(_06315_),
    .B1(_06338_),
    .C1(_06349_),
    .Y(_06351_));
 sky130_fd_sc_hd__o211ai_2 _12463_ (.A1(_06342_),
    .A2(_06346_),
    .B1(_06350_),
    .C1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__and2_1 _12464_ (.A(_06350_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__and2b_1 _12465_ (.A_N(_06353_),
    .B(_06314_),
    .X(_06354_));
 sky130_fd_sc_hd__a211o_1 _12466_ (.A1(_06350_),
    .A2(_06351_),
    .B1(_06342_),
    .C1(_06346_),
    .X(_06355_));
 sky130_fd_sc_hd__a2bb2o_1 _12467_ (.A1_N(_06346_),
    .A2_N(_06347_),
    .B1(_06348_),
    .B2(_06338_),
    .X(_06356_));
 sky130_fd_sc_hd__and2_1 _12468_ (.A(_06324_),
    .B(_06336_),
    .X(_06357_));
 sky130_fd_sc_hd__o2bb2a_1 _12469_ (.A1_N(net1611),
    .A2_N(net2239),
    .B1(_06318_),
    .B2(_06319_),
    .X(_06358_));
 sky130_fd_sc_hd__nor2_1 _12470_ (.A(_06320_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__and4_2 _12471_ (.A(net1607),
    .B(net1590),
    .C(net2078),
    .D(net2379),
    .X(_06360_));
 sky130_fd_sc_hd__a22o_1 _12472_ (.A1(net1607),
    .A2(net2078),
    .B1(net2379),
    .B2(net1590),
    .X(_06361_));
 sky130_fd_sc_hd__inv_2 _12473_ (.A(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__and4b_1 _12474_ (.A_N(_06360_),
    .B(_06361_),
    .C(net1632),
    .D(net821),
    .X(_06363_));
 sky130_fd_sc_hd__o2bb2a_1 _12475_ (.A1_N(net1632),
    .A2_N(net821),
    .B1(_06360_),
    .B2(_06362_),
    .X(_06364_));
 sky130_fd_sc_hd__nor2_1 _12476_ (.A(_06363_),
    .B(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_06359_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__nor3_1 _12478_ (.A(_06337_),
    .B(_06357_),
    .C(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__o21a_1 _12479_ (.A1(_06337_),
    .A2(_06357_),
    .B1(_06366_),
    .X(_06368_));
 sky130_fd_sc_hd__or2_1 _12480_ (.A(_06367_),
    .B(_06368_),
    .X(_06369_));
 sky130_fd_sc_hd__a22oi_1 _12481_ (.A1(net1574),
    .A2(net839),
    .B1(net2007),
    .B2(net1652),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _12482_ (.A(_04549_),
    .B(net2008),
    .Y(_06371_));
 sky130_fd_sc_hd__a22oi_1 _12483_ (.A1(net731),
    .A2(net1713),
    .B1(net1926),
    .B2(net914),
    .Y(_06372_));
 sky130_fd_sc_hd__nor2_1 _12484_ (.A(_04286_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__o21ai_2 _12485_ (.A1(_06360_),
    .A2(_06363_),
    .B1(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__or3_1 _12486_ (.A(_06360_),
    .B(_06363_),
    .C(_06373_),
    .X(_06375_));
 sky130_fd_sc_hd__and2_1 _12487_ (.A(_06374_),
    .B(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(net2009),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__or2_1 _12489_ (.A(net2009),
    .B(_06376_),
    .X(_06378_));
 sky130_fd_sc_hd__nand2_1 _12490_ (.A(net2010),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__nor2_1 _12491_ (.A(_06369_),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__o211a_1 _12492_ (.A1(_06367_),
    .A2(_06380_),
    .B1(_06349_),
    .C1(_06356_),
    .X(_06381_));
 sky130_fd_sc_hd__a211oi_1 _12493_ (.A1(_06349_),
    .A2(_06356_),
    .B1(_06367_),
    .C1(_06380_),
    .Y(_06382_));
 sky130_fd_sc_hd__or2_1 _12494_ (.A(_06381_),
    .B(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a21oi_1 _12495_ (.A1(_06374_),
    .A2(net2010),
    .B1(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__o211ai_2 _12496_ (.A1(_06381_),
    .A2(net2011),
    .B1(_06352_),
    .C1(_06355_),
    .Y(_06385_));
 sky130_fd_sc_hd__and3_1 _12497_ (.A(_06374_),
    .B(net2010),
    .C(_06383_),
    .X(_06386_));
 sky130_fd_sc_hd__and2_1 _12498_ (.A(_06369_),
    .B(_06379_),
    .X(_06387_));
 sky130_fd_sc_hd__nor2_1 _12499_ (.A(_06380_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__and4_2 _12500_ (.A(net1574),
    .B(net731),
    .C(net896),
    .D(net1926),
    .X(_06389_));
 sky130_fd_sc_hd__nand2_1 _12501_ (.A(_06388_),
    .B(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__or2_1 _12502_ (.A(_06359_),
    .B(_06365_),
    .X(_06391_));
 sky130_fd_sc_hd__nand2_1 _12503_ (.A(_06366_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__a22oi_2 _12504_ (.A1(net1574),
    .A2(net896),
    .B1(net1926),
    .B2(net731),
    .Y(_06393_));
 sky130_fd_sc_hd__nor3_1 _12505_ (.A(_06389_),
    .B(_06392_),
    .C(net3099),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _12506_ (.A(_06388_),
    .B(net3100),
    .Y(_06395_));
 sky130_fd_sc_hd__a211oi_2 _12507_ (.A1(_06390_),
    .A2(net3101),
    .B1(net2011),
    .C1(_06386_),
    .Y(_06396_));
 sky130_fd_sc_hd__a211o_1 _12508_ (.A1(_06352_),
    .A2(_06355_),
    .B1(_06381_),
    .C1(net2011),
    .X(_06397_));
 sky130_fd_sc_hd__nand3_1 _12509_ (.A(_06385_),
    .B(_06396_),
    .C(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__xor2_1 _12510_ (.A(_06314_),
    .B(_06353_),
    .X(_06399_));
 sky130_fd_sc_hd__a21oi_1 _12511_ (.A1(_06385_),
    .A2(_06398_),
    .B1(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__o21a_1 _12512_ (.A1(_06354_),
    .A2(_06400_),
    .B1(_06313_),
    .X(_06401_));
 sky130_fd_sc_hd__o21a_1 _12513_ (.A1(_06312_),
    .A2(_06401_),
    .B1(_06270_),
    .X(_06402_));
 sky130_fd_sc_hd__nor2_1 _12514_ (.A(_06268_),
    .B(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__xnor2_1 _12515_ (.A(_06230_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__xnor2_2 _12516_ (.A(_06228_),
    .B(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__o21ba_1 _12517_ (.A1(_06164_),
    .A2(_06174_),
    .B1_N(_06163_),
    .X(_06406_));
 sky130_fd_sc_hd__o21ai_1 _12518_ (.A1(_06117_),
    .A2(_06118_),
    .B1(_06121_),
    .Y(_06407_));
 sky130_fd_sc_hd__xnor2_1 _12519_ (.A(_06406_),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21oi_1 _12520_ (.A1(_06134_),
    .A2(_06136_),
    .B1(_06133_),
    .Y(_06409_));
 sky130_fd_sc_hd__a21o_1 _12521_ (.A1(_05462_),
    .A2(_05486_),
    .B1(_05458_),
    .X(_06410_));
 sky130_fd_sc_hd__xnor2_1 _12522_ (.A(_03518_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__xnor2_1 _12523_ (.A(_06409_),
    .B(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__xnor2_1 _12524_ (.A(_06408_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__and2b_1 _12525_ (.A_N(_03725_),
    .B(_03726_),
    .X(_06414_));
 sky130_fd_sc_hd__nand2b_1 _12526_ (.A_N(_05161_),
    .B(_05162_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_1 _12527_ (.A(_04889_),
    .B(_04928_),
    .Y(_06416_));
 sky130_fd_sc_hd__xnor2_1 _12528_ (.A(net3176),
    .B(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__xnor2_1 _12529_ (.A(_06414_),
    .B(net3177),
    .Y(_06418_));
 sky130_fd_sc_hd__xnor2_1 _12530_ (.A(_06413_),
    .B(net3178),
    .Y(_06419_));
 sky130_fd_sc_hd__xnor2_1 _12531_ (.A(_06405_),
    .B(net3179),
    .Y(_06420_));
 sky130_fd_sc_hd__xnor2_1 _12532_ (.A(net3678),
    .B(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(net1265),
    .A1(_06421_),
    .S(net37),
    .X(_00365_));
 sky130_fd_sc_hd__or3_1 _12534_ (.A(_06270_),
    .B(_06312_),
    .C(_06401_),
    .X(_06422_));
 sky130_fd_sc_hd__nor2_1 _12535_ (.A(net1247),
    .B(_06402_),
    .Y(_06423_));
 sky130_fd_sc_hd__a22o_1 _12536_ (.A1(net1151),
    .A2(net1247),
    .B1(_06422_),
    .B2(_06423_),
    .X(_00364_));
 sky130_fd_sc_hd__or3_1 _12537_ (.A(_06313_),
    .B(_06354_),
    .C(_06400_),
    .X(_06424_));
 sky130_fd_sc_hd__nor2_1 _12538_ (.A(net35),
    .B(_06401_),
    .Y(_06425_));
 sky130_fd_sc_hd__a22o_1 _12539_ (.A1(net299),
    .A2(net35),
    .B1(net2014),
    .B2(_06425_),
    .X(_00363_));
 sky130_fd_sc_hd__and3_1 _12540_ (.A(_06385_),
    .B(_06398_),
    .C(_06399_),
    .X(_06426_));
 sky130_fd_sc_hd__or2_1 _12541_ (.A(net35),
    .B(_06400_),
    .X(_06427_));
 sky130_fd_sc_hd__a2bb2o_1 _12542_ (.A1_N(_06426_),
    .A2_N(_06427_),
    .B1(net1259),
    .B2(net35),
    .X(_00362_));
 sky130_fd_sc_hd__and2_1 _12543_ (.A(net2552),
    .B(net35),
    .X(_06428_));
 sky130_fd_sc_hd__a21o_1 _12544_ (.A1(_06385_),
    .A2(_06397_),
    .B1(_06396_),
    .X(_06429_));
 sky130_fd_sc_hd__a31o_1 _12545_ (.A1(net250),
    .A2(net3103),
    .A3(_06429_),
    .B1(net2554),
    .X(_00361_));
 sky130_fd_sc_hd__o211a_1 _12546_ (.A1(net2011),
    .A2(_06386_),
    .B1(_06390_),
    .C1(_06395_),
    .X(_06430_));
 sky130_fd_sc_hd__or3_1 _12547_ (.A(net35),
    .B(_06396_),
    .C(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__a21bo_1 _12548_ (.A1(net1237),
    .A2(net35),
    .B1_N(_06431_),
    .X(_00360_));
 sky130_fd_sc_hd__or2_1 _12549_ (.A(_06388_),
    .B(_06394_),
    .X(_06432_));
 sky130_fd_sc_hd__and2_1 _12550_ (.A(_06395_),
    .B(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__o211a_1 _12551_ (.A1(_06389_),
    .A2(_06433_),
    .B1(_06390_),
    .C1(net250),
    .X(_06434_));
 sky130_fd_sc_hd__a21o_1 _12552_ (.A1(net1221),
    .A2(net35),
    .B1(_06434_),
    .X(_00359_));
 sky130_fd_sc_hd__o21a_1 _12553_ (.A1(_06389_),
    .A2(_06393_),
    .B1(_06392_),
    .X(_06435_));
 sky130_fd_sc_hd__or2_1 _12554_ (.A(net35),
    .B(_06394_),
    .X(_06436_));
 sky130_fd_sc_hd__a2bb2o_1 _12555_ (.A1_N(_06435_),
    .A2_N(_06436_),
    .B1(net1255),
    .B2(net35),
    .X(_00358_));
 sky130_fd_sc_hd__and2_2 _12556_ (.A(net1114),
    .B(net2634),
    .X(_06437_));
 sky130_fd_sc_hd__nand2_1 _12557_ (.A(net1114),
    .B(net2634),
    .Y(_06438_));
 sky130_fd_sc_hd__and3_1 _12558_ (.A(net2622),
    .B(net1110),
    .C(net2635),
    .X(_06439_));
 sky130_fd_sc_hd__nor2_1 _12559_ (.A(net1245),
    .B(net1110),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _12560_ (.A(net250),
    .B(net2636),
    .Y(_06441_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(net2636),
    .A1(_06441_),
    .S(net1184),
    .X(_00354_));
 sky130_fd_sc_hd__nor2_1 _12562_ (.A(net2622),
    .B(_06438_),
    .Y(_06442_));
 sky130_fd_sc_hd__a22o_1 _12563_ (.A1(net2622),
    .A2(_06441_),
    .B1(_06442_),
    .B2(net1110),
    .X(_00353_));
 sky130_fd_sc_hd__nor2_2 _12564_ (.A(net1114),
    .B(net2634),
    .Y(_06443_));
 sky130_fd_sc_hd__or2_4 _12565_ (.A(net1114),
    .B(net2634),
    .X(_06444_));
 sky130_fd_sc_hd__a32o_1 _12566_ (.A1(net1110),
    .A2(_06438_),
    .A3(_06444_),
    .B1(_06440_),
    .B2(net1114),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(net1110),
    .A1(_06440_),
    .S(net2634),
    .X(_00351_));
 sky130_fd_sc_hd__a21o_1 _12568_ (.A1(net1245),
    .A2(net1180),
    .B1(net1110),
    .X(_00350_));
 sky130_fd_sc_hd__a221o_1 _12569_ (.A1(net1289),
    .A2(_00668_),
    .B1(_06437_),
    .B2(net1233),
    .C1(_06443_),
    .X(_06445_));
 sky130_fd_sc_hd__and3b_1 _12570_ (.A_N(net2634),
    .B(net1114),
    .C(net1229),
    .X(_06446_));
 sky130_fd_sc_hd__o22a_1 _12571_ (.A1(net1138),
    .A2(_06444_),
    .B1(_06445_),
    .B2(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(net2646),
    .A1(net1139),
    .S(net1110),
    .X(_00349_));
 sky130_fd_sc_hd__a221o_1 _12573_ (.A1(net1285),
    .A2(_00668_),
    .B1(_06437_),
    .B2(net1321),
    .C1(_06443_),
    .X(_06448_));
 sky130_fd_sc_hd__and3b_1 _12574_ (.A_N(net2634),
    .B(net1114),
    .C(net1273),
    .X(_06449_));
 sky130_fd_sc_hd__o22a_1 _12575_ (.A1(net1151),
    .A2(_06444_),
    .B1(_06448_),
    .B2(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(net2651),
    .A1(net1152),
    .S(net1110),
    .X(_00348_));
 sky130_fd_sc_hd__a221o_1 _12577_ (.A1(net1269),
    .A2(_00668_),
    .B1(_06437_),
    .B2(net1325),
    .C1(_06443_),
    .X(_06451_));
 sky130_fd_sc_hd__and3b_1 _12578_ (.A_N(net2634),
    .B(net1114),
    .C(net1293),
    .X(_06452_));
 sky130_fd_sc_hd__o22a_1 _12579_ (.A1(net299),
    .A2(_06444_),
    .B1(_06451_),
    .B2(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(net2641),
    .A1(net296),
    .S(net1110),
    .X(_00347_));
 sky130_fd_sc_hd__a221o_1 _12581_ (.A1(net1251),
    .A2(_00668_),
    .B1(net2635),
    .B2(net2594),
    .C1(_06443_),
    .X(_06454_));
 sky130_fd_sc_hd__and3b_1 _12582_ (.A_N(net2634),
    .B(net1114),
    .C(net2564),
    .X(_06455_));
 sky130_fd_sc_hd__o22a_1 _12583_ (.A1(net1259),
    .A2(_06444_),
    .B1(_06454_),
    .B2(_06455_),
    .X(_06456_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(net1143),
    .A1(_06456_),
    .S(net1110),
    .X(_00346_));
 sky130_fd_sc_hd__a221o_1 _12585_ (.A1(net1415),
    .A2(_00668_),
    .B1(_06437_),
    .B2(net1317),
    .C1(_06443_),
    .X(_06457_));
 sky130_fd_sc_hd__and3b_1 _12586_ (.A_N(net704),
    .B(net1114),
    .C(net1313),
    .X(_06458_));
 sky130_fd_sc_hd__o22a_1 _12587_ (.A1(net2552),
    .A2(_06444_),
    .B1(_06457_),
    .B2(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(net2628),
    .A1(_06459_),
    .S(net1110),
    .X(_00345_));
 sky130_fd_sc_hd__a221o_1 _12589_ (.A1(net1211),
    .A2(_00668_),
    .B1(net2635),
    .B2(net1301),
    .C1(_06443_),
    .X(_06460_));
 sky130_fd_sc_hd__and3b_1 _12590_ (.A_N(net2634),
    .B(net1114),
    .C(net1305),
    .X(_06461_));
 sky130_fd_sc_hd__o22a_1 _12591_ (.A1(net1237),
    .A2(_06444_),
    .B1(_06460_),
    .B2(_06461_),
    .X(_06462_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(net1130),
    .A1(_06462_),
    .S(net1110),
    .X(_00344_));
 sky130_fd_sc_hd__a221o_1 _12593_ (.A1(net1225),
    .A2(_00668_),
    .B1(net2635),
    .B2(net2570),
    .C1(_06443_),
    .X(_06463_));
 sky130_fd_sc_hd__and3b_1 _12594_ (.A_N(net2634),
    .B(net1114),
    .C(net2546),
    .X(_06464_));
 sky130_fd_sc_hd__o22a_1 _12595_ (.A1(net1221),
    .A2(_06444_),
    .B1(_06463_),
    .B2(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(net1126),
    .A1(_06465_),
    .S(net1110),
    .X(_00343_));
 sky130_fd_sc_hd__mux4_2 _12597_ (.A0(net1255),
    .A1(net1188),
    .A2(net2558),
    .A3(net1397),
    .S0(net2634),
    .S1(net1114),
    .X(_06466_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(net1134),
    .A1(_06466_),
    .S(net1110),
    .X(_00342_));
 sky130_fd_sc_hd__nand2_4 _12599_ (.A(_03251_),
    .B(_03258_),
    .Y(_06467_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(net2368),
    .A1(net1999),
    .S(_06467_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(net1875),
    .A1(net2164),
    .S(_06467_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(net2327),
    .A1(net1942),
    .S(_06467_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(net1682),
    .A1(net2128),
    .S(_06467_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(net2033),
    .A1(net2119),
    .S(_06467_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(net2087),
    .A1(net2195),
    .S(_06467_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(net1797),
    .A1(net2045),
    .S(_06467_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(net1922),
    .A1(net2097),
    .S(_06467_),
    .X(_00334_));
 sky130_fd_sc_hd__or2_1 _12608_ (.A(net1207),
    .B(net250),
    .X(_00333_));
 sky130_fd_sc_hd__a31o_1 _12609_ (.A1(net19),
    .A2(_03243_),
    .A3(_03258_),
    .B1(_03264_),
    .X(_06468_));
 sky130_fd_sc_hd__or4_1 _12610_ (.A(net360),
    .B(net1198),
    .C(net1021),
    .D(net20),
    .X(_06469_));
 sky130_fd_sc_hd__a41o_1 _12611_ (.A1(net10),
    .A2(net1192),
    .A3(net1401),
    .A4(net1622),
    .B1(net1023),
    .X(_06470_));
 sky130_fd_sc_hd__and4_1 _12612_ (.A(_00000_),
    .B(_06468_),
    .C(_06469_),
    .D(net1193),
    .X(_06471_));
 sky130_fd_sc_hd__a21o_1 _12613_ (.A1(net1596),
    .A2(net1022),
    .B1(net360),
    .X(_06472_));
 sky130_fd_sc_hd__o211a_1 _12614_ (.A1(net1596),
    .A2(net1022),
    .B1(net1194),
    .C1(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__o21ba_1 _12615_ (.A1(net1217),
    .A2(net1194),
    .B1_N(net255),
    .X(_00355_));
 sky130_fd_sc_hd__xor2_1 _12616_ (.A(net1198),
    .B(net1021),
    .X(_06474_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(net1077),
    .A1(net244),
    .S(net1194),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _12618_ (.A0(net1199),
    .A1(net244),
    .S(net360),
    .X(_06475_));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(net1075),
    .A1(net1201),
    .S(net1194),
    .X(_00357_));
 sky130_fd_sc_hd__inv_2 _12620_ (.A(net198),
    .Y(_00001_));
 sky130_fd_sc_hd__inv_2 _12621_ (.A(net198),
    .Y(_00002_));
 sky130_fd_sc_hd__inv_2 _12622_ (.A(net196),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_2 _12623_ (.A(net191),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _12624_ (.A(net191),
    .Y(_00005_));
 sky130_fd_sc_hd__inv_2 _12625_ (.A(net191),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _12626_ (.A(net191),
    .Y(_00007_));
 sky130_fd_sc_hd__inv_2 _12627_ (.A(net191),
    .Y(_00008_));
 sky130_fd_sc_hd__inv_2 _12628_ (.A(net191),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _12629_ (.A(net191),
    .Y(_00010_));
 sky130_fd_sc_hd__inv_2 _12630_ (.A(net191),
    .Y(_00011_));
 sky130_fd_sc_hd__inv_2 _12631_ (.A(net202),
    .Y(_00012_));
 sky130_fd_sc_hd__inv_2 _12632_ (.A(net202),
    .Y(_00013_));
 sky130_fd_sc_hd__inv_2 _12633_ (.A(net196),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _12634_ (.A(net196),
    .Y(_00015_));
 sky130_fd_sc_hd__inv_2 _12635_ (.A(net196),
    .Y(_00016_));
 sky130_fd_sc_hd__inv_2 _12636_ (.A(net196),
    .Y(_00017_));
 sky130_fd_sc_hd__inv_2 _12637_ (.A(net209),
    .Y(_00018_));
 sky130_fd_sc_hd__inv_2 _12638_ (.A(net209),
    .Y(_00019_));
 sky130_fd_sc_hd__inv_2 _12639_ (.A(net202),
    .Y(_00020_));
 sky130_fd_sc_hd__inv_2 _12640_ (.A(net199),
    .Y(_00021_));
 sky130_fd_sc_hd__inv_2 _12641_ (.A(net199),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_2 _12642_ (.A(net199),
    .Y(_00023_));
 sky130_fd_sc_hd__inv_2 _12643_ (.A(net199),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_2 _12644_ (.A(net201),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_2 _12645_ (.A(net201),
    .Y(_00026_));
 sky130_fd_sc_hd__inv_2 _12646_ (.A(net199),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _12647_ (.A(net199),
    .Y(_00028_));
 sky130_fd_sc_hd__inv_2 _12648_ (.A(net199),
    .Y(_00029_));
 sky130_fd_sc_hd__inv_2 _12649_ (.A(net206),
    .Y(_00030_));
 sky130_fd_sc_hd__inv_2 _12650_ (.A(net209),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _12651_ (.A(net209),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_2 _12652_ (.A(net189),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_2 _12653_ (.A(net189),
    .Y(_00034_));
 sky130_fd_sc_hd__inv_2 _12654_ (.A(net189),
    .Y(_00035_));
 sky130_fd_sc_hd__inv_2 _12655_ (.A(net189),
    .Y(_00036_));
 sky130_fd_sc_hd__inv_2 _12656_ (.A(net189),
    .Y(_00037_));
 sky130_fd_sc_hd__inv_2 _12657_ (.A(net193),
    .Y(_00038_));
 sky130_fd_sc_hd__inv_2 _12658_ (.A(net193),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _12659_ (.A(net193),
    .Y(_00040_));
 sky130_fd_sc_hd__inv_2 _12660_ (.A(net201),
    .Y(_00041_));
 sky130_fd_sc_hd__inv_2 _12661_ (.A(net201),
    .Y(_00042_));
 sky130_fd_sc_hd__inv_2 _12662_ (.A(net201),
    .Y(_00043_));
 sky130_fd_sc_hd__inv_2 _12663_ (.A(net201),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_2 _12664_ (.A(net201),
    .Y(_00045_));
 sky130_fd_sc_hd__inv_2 _12665_ (.A(net209),
    .Y(_00046_));
 sky130_fd_sc_hd__inv_2 _12666_ (.A(net209),
    .Y(_00047_));
 sky130_fd_sc_hd__inv_2 _12667_ (.A(net209),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_2 _12668_ (.A(net203),
    .Y(_00049_));
 sky130_fd_sc_hd__inv_2 _12669_ (.A(net203),
    .Y(_00050_));
 sky130_fd_sc_hd__inv_2 _12670_ (.A(net203),
    .Y(_00051_));
 sky130_fd_sc_hd__inv_2 _12671_ (.A(net203),
    .Y(_00052_));
 sky130_fd_sc_hd__inv_2 _12672_ (.A(net196),
    .Y(_00053_));
 sky130_fd_sc_hd__inv_2 _12673_ (.A(net200),
    .Y(_00054_));
 sky130_fd_sc_hd__inv_2 _12674_ (.A(net202),
    .Y(_00055_));
 sky130_fd_sc_hd__inv_2 _12675_ (.A(net202),
    .Y(_00056_));
 sky130_fd_sc_hd__inv_2 _12676_ (.A(net208),
    .Y(_00057_));
 sky130_fd_sc_hd__inv_2 _12677_ (.A(net208),
    .Y(_00058_));
 sky130_fd_sc_hd__inv_2 _12678_ (.A(net208),
    .Y(_00059_));
 sky130_fd_sc_hd__inv_2 _12679_ (.A(net205),
    .Y(_00060_));
 sky130_fd_sc_hd__inv_2 _12680_ (.A(net194),
    .Y(_00061_));
 sky130_fd_sc_hd__inv_2 _12681_ (.A(net193),
    .Y(_00062_));
 sky130_fd_sc_hd__inv_2 _12682_ (.A(net193),
    .Y(_00063_));
 sky130_fd_sc_hd__inv_2 _12683_ (.A(net193),
    .Y(_00064_));
 sky130_fd_sc_hd__inv_2 _12684_ (.A(net203),
    .Y(_00065_));
 sky130_fd_sc_hd__inv_2 _12685_ (.A(net192),
    .Y(_00066_));
 sky130_fd_sc_hd__inv_2 _12686_ (.A(net192),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _12687_ (.A(net192),
    .Y(_00068_));
 sky130_fd_sc_hd__inv_2 _12688_ (.A(net192),
    .Y(_00069_));
 sky130_fd_sc_hd__inv_2 _12689_ (.A(net192),
    .Y(_00070_));
 sky130_fd_sc_hd__inv_2 _12690_ (.A(net191),
    .Y(_00071_));
 sky130_fd_sc_hd__inv_2 _12691_ (.A(net187),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_2 _12692_ (.A(net188),
    .Y(_00073_));
 sky130_fd_sc_hd__inv_2 _12693_ (.A(net203),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_2 _12694_ (.A(net193),
    .Y(_00075_));
 sky130_fd_sc_hd__inv_2 _12695_ (.A(net198),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _12696_ (.A(net194),
    .Y(_00077_));
 sky130_fd_sc_hd__inv_2 _12697_ (.A(net194),
    .Y(_00078_));
 sky130_fd_sc_hd__inv_2 _12698_ (.A(net194),
    .Y(_00079_));
 sky130_fd_sc_hd__inv_2 _12699_ (.A(net194),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _12700_ (.A(net194),
    .Y(_00081_));
 sky130_fd_sc_hd__inv_2 _12701_ (.A(net194),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _12702_ (.A(net194),
    .Y(_00083_));
 sky130_fd_sc_hd__inv_2 _12703_ (.A(net194),
    .Y(_00084_));
 sky130_fd_sc_hd__inv_2 _12704_ (.A(net194),
    .Y(_00085_));
 sky130_fd_sc_hd__inv_2 _12705_ (.A(net194),
    .Y(_00086_));
 sky130_fd_sc_hd__inv_2 _12706_ (.A(net194),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _12707_ (.A(net203),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_2 _12708_ (.A(net203),
    .Y(_00089_));
 sky130_fd_sc_hd__inv_2 _12709_ (.A(net203),
    .Y(_00090_));
 sky130_fd_sc_hd__inv_2 _12710_ (.A(net203),
    .Y(_00091_));
 sky130_fd_sc_hd__inv_2 _12711_ (.A(net205),
    .Y(_00092_));
 sky130_fd_sc_hd__inv_2 _12712_ (.A(net187),
    .Y(_00093_));
 sky130_fd_sc_hd__inv_2 _12713_ (.A(net187),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _12714_ (.A(net187),
    .Y(_00095_));
 sky130_fd_sc_hd__inv_2 _12715_ (.A(net187),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _12716_ (.A(net187),
    .Y(_00097_));
 sky130_fd_sc_hd__inv_2 _12717_ (.A(net187),
    .Y(_00098_));
 sky130_fd_sc_hd__inv_2 _12718_ (.A(net187),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_2 _12719_ (.A(net187),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _12720_ (.A(net193),
    .Y(_00101_));
 sky130_fd_sc_hd__inv_2 _12721_ (.A(net193),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _12722_ (.A(net191),
    .Y(_00103_));
 sky130_fd_sc_hd__inv_2 _12723_ (.A(net191),
    .Y(_00104_));
 sky130_fd_sc_hd__inv_2 _12724_ (.A(net191),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _12725_ (.A(net191),
    .Y(_00106_));
 sky130_fd_sc_hd__inv_2 _12726_ (.A(net191),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _12727_ (.A(net191),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _12728_ (.A(net187),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _12729_ (.A(net187),
    .Y(_00110_));
 sky130_fd_sc_hd__inv_2 _12730_ (.A(net187),
    .Y(_00111_));
 sky130_fd_sc_hd__inv_2 _12731_ (.A(net188),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_2 _12732_ (.A(net188),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _12733_ (.A(net188),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_2 _12734_ (.A(net188),
    .Y(_00115_));
 sky130_fd_sc_hd__inv_2 _12735_ (.A(net188),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_2 _12736_ (.A(net198),
    .Y(_00117_));
 sky130_fd_sc_hd__inv_2 _12737_ (.A(net198),
    .Y(_00118_));
 sky130_fd_sc_hd__inv_2 _12738_ (.A(net198),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _12739_ (.A(net197),
    .Y(_00120_));
 sky130_fd_sc_hd__inv_2 _12740_ (.A(net197),
    .Y(_00121_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(net198),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _12742_ (.A(net197),
    .Y(_00123_));
 sky130_fd_sc_hd__inv_2 _12743_ (.A(net197),
    .Y(_00124_));
 sky130_fd_sc_hd__inv_2 _12744_ (.A(net189),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _12745_ (.A(net189),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _12746_ (.A(net189),
    .Y(_00127_));
 sky130_fd_sc_hd__inv_2 _12747_ (.A(net190),
    .Y(_00128_));
 sky130_fd_sc_hd__inv_2 _12748_ (.A(net190),
    .Y(_00129_));
 sky130_fd_sc_hd__inv_2 _12749_ (.A(net190),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_2 _12750_ (.A(net190),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _12751_ (.A(net190),
    .Y(_00132_));
 sky130_fd_sc_hd__inv_2 _12752_ (.A(net208),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_2 _12753_ (.A(net208),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _12754_ (.A(net208),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _12755_ (.A(net207),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_2 _12756_ (.A(net207),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_2 _12757_ (.A(net207),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_2 _12758_ (.A(net207),
    .Y(_00139_));
 sky130_fd_sc_hd__inv_2 _12759_ (.A(net208),
    .Y(_00140_));
 sky130_fd_sc_hd__inv_2 _12760_ (.A(net205),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _12761_ (.A(net205),
    .Y(_00142_));
 sky130_fd_sc_hd__inv_2 _12762_ (.A(net205),
    .Y(_00143_));
 sky130_fd_sc_hd__inv_2 _12763_ (.A(net205),
    .Y(_00144_));
 sky130_fd_sc_hd__inv_2 _12764_ (.A(net205),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _12765_ (.A(net205),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _12766_ (.A(net205),
    .Y(_00147_));
 sky130_fd_sc_hd__inv_2 _12767_ (.A(net205),
    .Y(_00148_));
 sky130_fd_sc_hd__inv_2 _12768_ (.A(net209),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _12769_ (.A(net209),
    .Y(_00150_));
 sky130_fd_sc_hd__inv_2 _12770_ (.A(net207),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _12771_ (.A(net207),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _12772_ (.A(net207),
    .Y(_00153_));
 sky130_fd_sc_hd__inv_2 _12773_ (.A(net207),
    .Y(_00154_));
 sky130_fd_sc_hd__inv_2 _12774_ (.A(net207),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _12775_ (.A(net207),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _12776_ (.A(net198),
    .Y(_00157_));
 sky130_fd_sc_hd__inv_2 _12777_ (.A(net198),
    .Y(_00158_));
 sky130_fd_sc_hd__inv_2 _12778_ (.A(net198),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _12779_ (.A(net198),
    .Y(_00160_));
 sky130_fd_sc_hd__inv_2 _12780_ (.A(net198),
    .Y(_00161_));
 sky130_fd_sc_hd__inv_2 _12781_ (.A(net197),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _12782_ (.A(net197),
    .Y(_00163_));
 sky130_fd_sc_hd__inv_2 _12783_ (.A(net197),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _12784_ (.A(net203),
    .Y(_00165_));
 sky130_fd_sc_hd__inv_2 _12785_ (.A(net203),
    .Y(_00166_));
 sky130_fd_sc_hd__inv_2 _12786_ (.A(net203),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _12787_ (.A(net204),
    .Y(_00168_));
 sky130_fd_sc_hd__inv_2 _12788_ (.A(net204),
    .Y(_00169_));
 sky130_fd_sc_hd__inv_2 _12789_ (.A(net204),
    .Y(_00170_));
 sky130_fd_sc_hd__inv_2 _12790_ (.A(net204),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _12791_ (.A(net204),
    .Y(_00172_));
 sky130_fd_sc_hd__inv_2 _12792_ (.A(net201),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _12793_ (.A(net200),
    .Y(_00174_));
 sky130_fd_sc_hd__inv_2 _12794_ (.A(net200),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _12795_ (.A(net200),
    .Y(_00176_));
 sky130_fd_sc_hd__inv_2 _12796_ (.A(net200),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _12797_ (.A(net200),
    .Y(_00178_));
 sky130_fd_sc_hd__inv_2 _12798_ (.A(net200),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _12799_ (.A(net200),
    .Y(_00180_));
 sky130_fd_sc_hd__inv_2 _12800_ (.A(net199),
    .Y(_00181_));
 sky130_fd_sc_hd__inv_2 _12801_ (.A(net201),
    .Y(_00182_));
 sky130_fd_sc_hd__inv_2 _12802_ (.A(net201),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _12803_ (.A(net201),
    .Y(_00184_));
 sky130_fd_sc_hd__inv_2 _12804_ (.A(net202),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _12805_ (.A(net202),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _12806_ (.A(net202),
    .Y(_00187_));
 sky130_fd_sc_hd__inv_2 _12807_ (.A(net202),
    .Y(_00188_));
 sky130_fd_sc_hd__inv_2 _12808_ (.A(net199),
    .Y(_00189_));
 sky130_fd_sc_hd__inv_2 _12809_ (.A(net199),
    .Y(_00190_));
 sky130_fd_sc_hd__inv_2 _12810_ (.A(net199),
    .Y(_00191_));
 sky130_fd_sc_hd__inv_2 _12811_ (.A(net196),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _12812_ (.A(net196),
    .Y(_00193_));
 sky130_fd_sc_hd__inv_2 _12813_ (.A(net196),
    .Y(_00194_));
 sky130_fd_sc_hd__inv_2 _12814_ (.A(net196),
    .Y(_00195_));
 sky130_fd_sc_hd__inv_2 _12815_ (.A(net196),
    .Y(_00196_));
 sky130_fd_sc_hd__inv_2 _12816_ (.A(net193),
    .Y(_00197_));
 sky130_fd_sc_hd__inv_2 _12817_ (.A(net193),
    .Y(_00198_));
 sky130_fd_sc_hd__inv_2 _12818_ (.A(net193),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _12819_ (.A(net193),
    .Y(_00200_));
 sky130_fd_sc_hd__inv_2 _12820_ (.A(net192),
    .Y(_00201_));
 sky130_fd_sc_hd__inv_2 _12821_ (.A(net192),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _12822_ (.A(net192),
    .Y(_00203_));
 sky130_fd_sc_hd__inv_2 _12823_ (.A(net192),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _12824_ (.A(net189),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _12825_ (.A(net189),
    .Y(_00206_));
 sky130_fd_sc_hd__inv_2 _12826_ (.A(net195),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _12827_ (.A(net195),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_2 _12828_ (.A(net189),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _12829_ (.A(net189),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _12830_ (.A(net189),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _12831_ (.A(net195),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _12832_ (.A(net194),
    .Y(_00213_));
 sky130_fd_sc_hd__inv_2 _12833_ (.A(net194),
    .Y(_00214_));
 sky130_fd_sc_hd__inv_2 _12834_ (.A(net194),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _12835_ (.A(net195),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _12836_ (.A(net195),
    .Y(_00217_));
 sky130_fd_sc_hd__inv_2 _12837_ (.A(net195),
    .Y(_00218_));
 sky130_fd_sc_hd__inv_2 _12838_ (.A(net195),
    .Y(_00219_));
 sky130_fd_sc_hd__inv_2 _12839_ (.A(net195),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _12840_ (.A(net204),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _12841_ (.A(net204),
    .Y(_00222_));
 sky130_fd_sc_hd__inv_2 _12842_ (.A(net204),
    .Y(_00223_));
 sky130_fd_sc_hd__inv_2 _12843_ (.A(net203),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _12844_ (.A(net204),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_2 _12845_ (.A(net204),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _12846_ (.A(net204),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _12847_ (.A(net204),
    .Y(_00228_));
 sky130_fd_sc_hd__inv_2 _12848_ (.A(net189),
    .Y(_00229_));
 sky130_fd_sc_hd__inv_2 _12849_ (.A(net189),
    .Y(_00230_));
 sky130_fd_sc_hd__inv_2 _12850_ (.A(net187),
    .Y(_00231_));
 sky130_fd_sc_hd__inv_2 _12851_ (.A(net187),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _12852_ (.A(net187),
    .Y(_00233_));
 sky130_fd_sc_hd__inv_2 _12853_ (.A(net187),
    .Y(_00234_));
 sky130_fd_sc_hd__inv_2 _12854_ (.A(net188),
    .Y(_00235_));
 sky130_fd_sc_hd__inv_2 _12855_ (.A(net188),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _12856_ (.A(net193),
    .Y(_00237_));
 sky130_fd_sc_hd__inv_2 _12857_ (.A(net193),
    .Y(_00238_));
 sky130_fd_sc_hd__inv_2 _12858_ (.A(net193),
    .Y(_00239_));
 sky130_fd_sc_hd__inv_2 _12859_ (.A(net191),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _12860_ (.A(net192),
    .Y(_00241_));
 sky130_fd_sc_hd__inv_2 _12861_ (.A(net192),
    .Y(_00242_));
 sky130_fd_sc_hd__inv_2 _12862_ (.A(net192),
    .Y(_00243_));
 sky130_fd_sc_hd__inv_2 _12863_ (.A(net192),
    .Y(_00244_));
 sky130_fd_sc_hd__inv_2 _12864_ (.A(net189),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _12865_ (.A(net190),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _12866_ (.A(net188),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _12867_ (.A(net188),
    .Y(_00248_));
 sky130_fd_sc_hd__inv_2 _12868_ (.A(net188),
    .Y(_00249_));
 sky130_fd_sc_hd__inv_2 _12869_ (.A(net190),
    .Y(_00250_));
 sky130_fd_sc_hd__inv_2 _12870_ (.A(net190),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _12871_ (.A(net188),
    .Y(_00252_));
 sky130_fd_sc_hd__inv_2 _12872_ (.A(net199),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_2 _12873_ (.A(net197),
    .Y(_00254_));
 sky130_fd_sc_hd__inv_2 _12874_ (.A(net197),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_2 _12875_ (.A(net197),
    .Y(_00256_));
 sky130_fd_sc_hd__inv_2 _12876_ (.A(net197),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _12877_ (.A(net197),
    .Y(_00258_));
 sky130_fd_sc_hd__inv_2 _12878_ (.A(net197),
    .Y(_00259_));
 sky130_fd_sc_hd__inv_2 _12879_ (.A(net197),
    .Y(_00260_));
 sky130_fd_sc_hd__inv_2 _12880_ (.A(net195),
    .Y(_00261_));
 sky130_fd_sc_hd__inv_2 _12881_ (.A(net190),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _12882_ (.A(net190),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _12883_ (.A(net190),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _12884_ (.A(net190),
    .Y(_00265_));
 sky130_fd_sc_hd__inv_2 _12885_ (.A(net190),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _12886_ (.A(net190),
    .Y(_00267_));
 sky130_fd_sc_hd__inv_2 _12887_ (.A(net190),
    .Y(_00268_));
 sky130_fd_sc_hd__inv_2 _12888_ (.A(net209),
    .Y(_00269_));
 sky130_fd_sc_hd__inv_2 _12889_ (.A(net209),
    .Y(_00270_));
 sky130_fd_sc_hd__inv_2 _12890_ (.A(net208),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _12891_ (.A(net208),
    .Y(_00272_));
 sky130_fd_sc_hd__inv_2 _12892_ (.A(net208),
    .Y(_00273_));
 sky130_fd_sc_hd__inv_2 _12893_ (.A(net208),
    .Y(_00274_));
 sky130_fd_sc_hd__inv_2 _12894_ (.A(net208),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _12895_ (.A(net208),
    .Y(_00276_));
 sky130_fd_sc_hd__inv_2 _12896_ (.A(net206),
    .Y(_00277_));
 sky130_fd_sc_hd__inv_2 _12897_ (.A(net206),
    .Y(_00278_));
 sky130_fd_sc_hd__inv_2 _12898_ (.A(net205),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _12899_ (.A(net206),
    .Y(_00280_));
 sky130_fd_sc_hd__inv_2 _12900_ (.A(net206),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _12901_ (.A(net206),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _12902_ (.A(net206),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _12903_ (.A(net206),
    .Y(_00284_));
 sky130_fd_sc_hd__inv_2 _12904_ (.A(net209),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _12905_ (.A(net209),
    .Y(_00286_));
 sky130_fd_sc_hd__inv_2 _12906_ (.A(net207),
    .Y(_00287_));
 sky130_fd_sc_hd__inv_2 _12907_ (.A(net207),
    .Y(_00288_));
 sky130_fd_sc_hd__inv_2 _12908_ (.A(net207),
    .Y(_00289_));
 sky130_fd_sc_hd__inv_2 _12909_ (.A(net207),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _12910_ (.A(net207),
    .Y(_00291_));
 sky130_fd_sc_hd__inv_2 _12911_ (.A(net207),
    .Y(_00292_));
 sky130_fd_sc_hd__inv_2 _12912_ (.A(net198),
    .Y(_00293_));
 sky130_fd_sc_hd__inv_2 _12913_ (.A(net198),
    .Y(_00294_));
 sky130_fd_sc_hd__inv_2 _12914_ (.A(net198),
    .Y(_00295_));
 sky130_fd_sc_hd__inv_2 _12915_ (.A(net198),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _12916_ (.A(net197),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _12917_ (.A(net197),
    .Y(_00298_));
 sky130_fd_sc_hd__inv_2 _12918_ (.A(net210),
    .Y(_00299_));
 sky130_fd_sc_hd__inv_2 _12919_ (.A(net210),
    .Y(_00300_));
 sky130_fd_sc_hd__inv_2 _12920_ (.A(net203),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _12921_ (.A(net204),
    .Y(_00302_));
 sky130_fd_sc_hd__inv_2 _12922_ (.A(net204),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _12923_ (.A(net205),
    .Y(_00304_));
 sky130_fd_sc_hd__inv_2 _12924_ (.A(net205),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _12925_ (.A(net205),
    .Y(_00306_));
 sky130_fd_sc_hd__inv_2 _12926_ (.A(net205),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _12927_ (.A(net205),
    .Y(_00308_));
 sky130_fd_sc_hd__inv_2 _12928_ (.A(net200),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _12929_ (.A(net200),
    .Y(_00310_));
 sky130_fd_sc_hd__inv_2 _12930_ (.A(net200),
    .Y(_00311_));
 sky130_fd_sc_hd__inv_2 _12931_ (.A(net200),
    .Y(_00312_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(net200),
    .Y(_00313_));
 sky130_fd_sc_hd__inv_2 _12933_ (.A(net200),
    .Y(_00314_));
 sky130_fd_sc_hd__inv_2 _12934_ (.A(net201),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _12935_ (.A(net201),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _12936_ (.A(net199),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _12937_ (.A(net202),
    .Y(_00318_));
 sky130_fd_sc_hd__inv_2 _12938_ (.A(net202),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _12939_ (.A(net202),
    .Y(_00320_));
 sky130_fd_sc_hd__inv_2 _12940_ (.A(net202),
    .Y(_00321_));
 sky130_fd_sc_hd__inv_2 _12941_ (.A(net202),
    .Y(_00322_));
 sky130_fd_sc_hd__inv_2 _12942_ (.A(net200),
    .Y(_00323_));
 sky130_fd_sc_hd__inv_2 _12943_ (.A(net200),
    .Y(_00324_));
 sky130_fd_sc_hd__inv_2 _12944_ (.A(net199),
    .Y(_00325_));
 sky130_fd_sc_hd__inv_2 _12945_ (.A(net196),
    .Y(_00326_));
 sky130_fd_sc_hd__inv_2 _12946_ (.A(net196),
    .Y(_00327_));
 sky130_fd_sc_hd__inv_2 _12947_ (.A(net196),
    .Y(_00328_));
 sky130_fd_sc_hd__inv_2 _12948_ (.A(net196),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _12949_ (.A(net196),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_2 _12950_ (.A(net202),
    .Y(_00331_));
 sky130_fd_sc_hd__inv_2 _12951_ (.A(net202),
    .Y(_00332_));
 sky130_fd_sc_hd__dfrtp_1 _12952_ (.CLK(clknet_leaf_24_clk),
    .D(net1217),
    .RESET_B(_00000_),
    .Q(\control_fsm.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12953_ (.CLK(clknet_leaf_4_clk),
    .D(net2620),
    .RESET_B(_00001_),
    .Q(\control_fsm.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12954_ (.CLK(clknet_leaf_24_clk),
    .D(net2616),
    .RESET_B(_00002_),
    .Q(\control_fsm.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12955_ (.CLK(clknet_leaf_7_clk),
    .D(net1209),
    .RESET_B(_00003_),
    .Q(\next_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12956_ (.CLK(clknet_leaf_55_clk),
    .D(net2099),
    .RESET_B(_00004_),
    .Q(\mac_array.mac[15].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12957_ (.CLK(clknet_leaf_56_clk),
    .D(net2047),
    .RESET_B(_00005_),
    .Q(\mac_array.mac[15].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12958_ (.CLK(clknet_leaf_56_clk),
    .D(net2197),
    .RESET_B(_00006_),
    .Q(\mac_array.mac[15].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12959_ (.CLK(clknet_leaf_51_clk),
    .D(net2121),
    .RESET_B(_00007_),
    .Q(\mac_array.mac[15].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12960_ (.CLK(clknet_leaf_51_clk),
    .D(net2130),
    .RESET_B(_00008_),
    .Q(\mac_array.mac[15].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12961_ (.CLK(clknet_leaf_51_clk),
    .D(net1944),
    .RESET_B(_00009_),
    .Q(\mac_array.mac[15].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12962_ (.CLK(clknet_leaf_51_clk),
    .D(net2166),
    .RESET_B(_00010_),
    .Q(\mac_array.mac[15].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12963_ (.CLK(clknet_leaf_51_clk),
    .D(net2001),
    .RESET_B(_00011_),
    .Q(\mac_array.mac[15].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12964_ (.CLK(clknet_leaf_13_clk),
    .D(net1136),
    .RESET_B(_00012_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_4 _12965_ (.CLK(clknet_leaf_13_clk),
    .D(net1128),
    .RESET_B(_00013_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_4 _12966_ (.CLK(clknet_leaf_12_clk),
    .D(net1132),
    .RESET_B(_00014_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_4 _12967_ (.CLK(clknet_leaf_11_clk),
    .D(net2632),
    .RESET_B(_00015_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_4 _12968_ (.CLK(clknet_leaf_7_clk),
    .D(net1145),
    .RESET_B(_00016_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_4 _12969_ (.CLK(clknet_leaf_11_clk),
    .D(net1099),
    .RESET_B(_00017_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_4 _12970_ (.CLK(clknet_leaf_28_clk),
    .D(net1154),
    .RESET_B(_00018_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_4 _12971_ (.CLK(clknet_leaf_28_clk),
    .D(net1141),
    .RESET_B(_00019_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_4 _12972_ (.CLK(clknet_3_5__leaf_clk),
    .D(net1182),
    .RESET_B(_00020_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _12973_ (.CLK(clknet_leaf_23_clk),
    .D(net1112),
    .RESET_B(_00021_),
    .Q(\result_index[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12974_ (.CLK(clknet_leaf_23_clk),
    .D(net1116),
    .RESET_B(_00022_),
    .Q(\result_index[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12975_ (.CLK(clknet_leaf_23_clk),
    .D(net2626),
    .RESET_B(_00023_),
    .Q(\result_index[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12976_ (.CLK(clknet_leaf_22_clk),
    .D(net1186),
    .RESET_B(_00024_),
    .Q(\result_index[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_24_clk),
    .D(net1219),
    .Q(\control_fsm.next_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_4_clk),
    .D(net1196),
    .Q(\control_fsm.next_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_4_clk),
    .D(net1203),
    .Q(\control_fsm.next_state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12980_ (.CLK(clknet_leaf_22_clk),
    .D(net1257),
    .RESET_B(_00025_),
    .Q(\result[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _12981_ (.CLK(clknet_leaf_21_clk),
    .D(net1223),
    .RESET_B(_00026_),
    .Q(\result[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _12982_ (.CLK(clknet_leaf_23_clk),
    .D(net1239),
    .RESET_B(_00027_),
    .Q(\result[0][2] ));
 sky130_fd_sc_hd__dfrtp_1 _12983_ (.CLK(clknet_leaf_23_clk),
    .D(net2556),
    .RESET_B(_00028_),
    .Q(\result[0][3] ));
 sky130_fd_sc_hd__dfrtp_1 _12984_ (.CLK(clknet_leaf_23_clk),
    .D(net1261),
    .RESET_B(_00029_),
    .Q(\result[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _12985_ (.CLK(clknet_3_6__leaf_clk),
    .D(net2016),
    .RESET_B(_00030_),
    .Q(\result[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _12986_ (.CLK(clknet_leaf_28_clk),
    .D(net1249),
    .RESET_B(_00031_),
    .Q(\result[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _12987_ (.CLK(clknet_leaf_28_clk),
    .D(net1267),
    .RESET_B(_00032_),
    .Q(\result[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _12988_ (.CLK(clknet_leaf_3_clk),
    .D(net1190),
    .RESET_B(_00033_),
    .Q(\result[13][0] ));
 sky130_fd_sc_hd__dfrtp_1 _12989_ (.CLK(clknet_leaf_3_clk),
    .D(net1227),
    .RESET_B(_00034_),
    .Q(\result[13][1] ));
 sky130_fd_sc_hd__dfrtp_1 _12990_ (.CLK(clknet_leaf_4_clk),
    .D(net1213),
    .RESET_B(_00035_),
    .Q(\result[13][2] ));
 sky130_fd_sc_hd__dfrtp_1 _12991_ (.CLK(clknet_leaf_4_clk),
    .D(net1419),
    .RESET_B(_00036_),
    .Q(\result[13][3] ));
 sky130_fd_sc_hd__dfrtp_1 _12992_ (.CLK(clknet_leaf_59_clk),
    .D(net1253),
    .RESET_B(_00037_),
    .Q(\result[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _12993_ (.CLK(clknet_leaf_59_clk),
    .D(net1271),
    .RESET_B(_00038_),
    .Q(\result[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _12994_ (.CLK(clknet_leaf_59_clk),
    .D(net1287),
    .RESET_B(_00039_),
    .Q(\result[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _12995_ (.CLK(clknet_leaf_43_clk),
    .D(net1291),
    .RESET_B(_00040_),
    .Q(\result[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _12996_ (.CLK(clknet_leaf_21_clk),
    .D(net2562),
    .RESET_B(_00041_),
    .Q(\result[10][0] ));
 sky130_fd_sc_hd__dfrtp_1 _12997_ (.CLK(clknet_leaf_21_clk),
    .D(net2550),
    .RESET_B(_00042_),
    .Q(\result[10][1] ));
 sky130_fd_sc_hd__dfrtp_1 _12998_ (.CLK(clknet_leaf_21_clk),
    .D(net1307),
    .RESET_B(_00043_),
    .Q(\result[10][2] ));
 sky130_fd_sc_hd__dfrtp_1 _12999_ (.CLK(clknet_leaf_21_clk),
    .D(net1315),
    .RESET_B(_00044_),
    .Q(\result[10][3] ));
 sky130_fd_sc_hd__dfrtp_1 _13000_ (.CLK(clknet_leaf_21_clk),
    .D(net2568),
    .RESET_B(_00045_),
    .Q(\result[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _13001_ (.CLK(clknet_leaf_28_clk),
    .D(net1295),
    .RESET_B(_00046_),
    .Q(\result[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _13002_ (.CLK(clknet_leaf_28_clk),
    .D(net1275),
    .RESET_B(_00047_),
    .Q(\result[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _13003_ (.CLK(clknet_leaf_21_clk),
    .D(net1231),
    .RESET_B(_00048_),
    .Q(\result[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _13004_ (.CLK(clknet_leaf_42_clk),
    .D(net1446),
    .RESET_B(_00049_),
    .Q(\control_fsm.line_write_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13005_ (.CLK(clknet_leaf_42_clk),
    .D(net390),
    .RESET_B(_00050_),
    .Q(\control_fsm.line_write_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13006_ (.CLK(clknet_leaf_24_clk),
    .D(net1523),
    .RESET_B(_00051_),
    .Q(\control_fsm.line_write_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13007_ (.CLK(clknet_leaf_42_clk),
    .D(net1624),
    .RESET_B(_00052_),
    .Q(\control_fsm.line_write_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13008_ (.CLK(clknet_leaf_7_clk),
    .D(net1207),
    .RESET_B(_00053_),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13009_ (.CLK(clknet_leaf_18_clk),
    .D(net1375),
    .RESET_B(_00054_),
    .Q(\control_fsm.line_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13010_ (.CLK(clknet_leaf_15_clk),
    .D(net1566),
    .RESET_B(_00055_),
    .Q(\control_fsm.line_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13011_ (.CLK(clknet_leaf_15_clk),
    .D(net1556),
    .RESET_B(_00056_),
    .Q(\control_fsm.line_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13012_ (.CLK(clknet_leaf_33_clk),
    .D(net1019),
    .RESET_B(_00057_),
    .Q(\control_fsm.line_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13013_ (.CLK(clknet_leaf_33_clk),
    .D(net1015),
    .RESET_B(_00058_),
    .Q(\control_fsm.line_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13014_ (.CLK(clknet_leaf_33_clk),
    .D(net1025),
    .RESET_B(_00059_),
    .Q(\control_fsm.line_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13015_ (.CLK(clknet_3_6__leaf_clk),
    .D(net1391),
    .RESET_B(_00060_),
    .Q(\control_fsm.line_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13016_ (.CLK(clknet_3_3__leaf_clk),
    .D(net1379),
    .RESET_B(_00061_),
    .Q(\control_fsm.line_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13017_ (.CLK(clknet_leaf_43_clk),
    .D(net1896),
    .RESET_B(_00062_),
    .Q(\control_fsm.weight_write_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13018_ (.CLK(clknet_leaf_59_clk),
    .D(net1601),
    .RESET_B(_00063_),
    .Q(\control_fsm.weight_write_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13019_ (.CLK(clknet_leaf_43_clk),
    .D(net1548),
    .RESET_B(_00064_),
    .Q(\control_fsm.weight_write_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13020_ (.CLK(clknet_leaf_43_clk),
    .D(net1343),
    .RESET_B(_00065_),
    .Q(\control_fsm.weight_write_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13021_ (.CLK(clknet_leaf_50_clk),
    .D(net1073),
    .RESET_B(_00066_),
    .Q(\control_fsm.weight_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13022_ (.CLK(clknet_leaf_50_clk),
    .D(net1049),
    .RESET_B(_00067_),
    .Q(\control_fsm.weight_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13023_ (.CLK(clknet_leaf_50_clk),
    .D(net1043),
    .RESET_B(_00068_),
    .Q(\control_fsm.weight_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13024_ (.CLK(clknet_leaf_50_clk),
    .D(net1037),
    .RESET_B(_00069_),
    .Q(\control_fsm.weight_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13025_ (.CLK(clknet_3_2__leaf_clk),
    .D(net1055),
    .RESET_B(_00070_),
    .Q(\control_fsm.weight_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13026_ (.CLK(clknet_leaf_54_clk),
    .D(net1031),
    .RESET_B(_00071_),
    .Q(\control_fsm.weight_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13027_ (.CLK(clknet_3_0__leaf_clk),
    .D(net1061),
    .RESET_B(_00072_),
    .Q(\control_fsm.weight_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13028_ (.CLK(clknet_3_0__leaf_clk),
    .D(net1067),
    .RESET_B(_00073_),
    .Q(\control_fsm.weight_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13029_ (.CLK(clknet_leaf_24_clk),
    .D(net1339),
    .RESET_B(_00074_),
    .Q(\control_fsm.line_write_enable ));
 sky130_fd_sc_hd__dfrtp_1 _13030_ (.CLK(clknet_leaf_4_clk),
    .D(net1539),
    .RESET_B(_00075_),
    .Q(\control_fsm.weight_write_enable ));
 sky130_fd_sc_hd__dfrtp_4 _13031_ (.CLK(clknet_leaf_24_clk),
    .D(net1582),
    .RESET_B(_00076_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _13032_ (.CLK(clknet_leaf_46_clk),
    .D(net1727),
    .RESET_B(_00077_),
    .Q(\mac_array.mac[14].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13033_ (.CLK(clknet_leaf_46_clk),
    .D(net2108),
    .RESET_B(_00078_),
    .Q(\mac_array.mac[14].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13034_ (.CLK(clknet_leaf_46_clk),
    .D(net2089),
    .RESET_B(_00079_),
    .Q(\mac_array.mac[14].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13035_ (.CLK(clknet_leaf_46_clk),
    .D(net1835),
    .RESET_B(_00080_),
    .Q(\mac_array.mac[14].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13036_ (.CLK(clknet_leaf_44_clk),
    .D(net2093),
    .RESET_B(_00081_),
    .Q(\mac_array.mac[14].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13037_ (.CLK(clknet_leaf_46_clk),
    .D(net2125),
    .RESET_B(_00082_),
    .Q(\mac_array.mac[14].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13038_ (.CLK(clknet_leaf_46_clk),
    .D(net1919),
    .RESET_B(_00083_),
    .Q(\mac_array.mac[14].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13039_ (.CLK(clknet_leaf_46_clk),
    .D(net1355),
    .RESET_B(_00084_),
    .Q(\mac_array.mac[14].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13040_ (.CLK(clknet_leaf_43_clk),
    .D(net2146),
    .RESET_B(_00085_),
    .Q(\mac_array.mac[13].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13041_ (.CLK(clknet_leaf_43_clk),
    .D(net1090),
    .RESET_B(_00086_),
    .Q(\mac_array.mac[13].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13042_ (.CLK(clknet_leaf_43_clk),
    .D(net1084),
    .RESET_B(_00087_),
    .Q(\mac_array.mac[13].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13043_ (.CLK(clknet_leaf_42_clk),
    .D(net1178),
    .RESET_B(_00088_),
    .Q(\mac_array.mac[13].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13044_ (.CLK(clknet_leaf_42_clk),
    .D(net1684),
    .RESET_B(_00089_),
    .Q(\mac_array.mac[13].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13045_ (.CLK(clknet_leaf_41_clk),
    .D(net1087),
    .RESET_B(_00090_),
    .Q(\mac_array.mac[13].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13046_ (.CLK(clknet_leaf_41_clk),
    .D(net1166),
    .RESET_B(_00091_),
    .Q(\mac_array.mac[13].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13047_ (.CLK(clknet_leaf_41_clk),
    .D(net1093),
    .RESET_B(_00092_),
    .Q(\mac_array.mac[13].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13048_ (.CLK(clknet_leaf_61_clk),
    .D(net2043),
    .RESET_B(_00093_),
    .Q(\mac_array.mac[12].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13049_ (.CLK(clknet_leaf_62_clk),
    .D(net2544),
    .RESET_B(_00094_),
    .Q(\mac_array.mac[12].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13050_ (.CLK(clknet_leaf_62_clk),
    .D(net1731),
    .RESET_B(_00095_),
    .Q(\mac_array.mac[12].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13051_ (.CLK(clknet_leaf_62_clk),
    .D(net2532),
    .RESET_B(_00096_),
    .Q(\mac_array.mac[12].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13052_ (.CLK(clknet_leaf_62_clk),
    .D(net2526),
    .RESET_B(_00097_),
    .Q(\mac_array.mac[12].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13053_ (.CLK(clknet_leaf_62_clk),
    .D(net1843),
    .RESET_B(_00098_),
    .Q(\mac_array.mac[12].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13054_ (.CLK(clknet_leaf_62_clk),
    .D(net2417),
    .RESET_B(_00099_),
    .Q(\mac_array.mac[12].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13055_ (.CLK(clknet_leaf_62_clk),
    .D(net2509),
    .RESET_B(_00100_),
    .Q(\mac_array.mac[12].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13056_ (.CLK(clknet_leaf_58_clk),
    .D(net1915),
    .RESET_B(_00101_),
    .Q(\mac_array.mac[11].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13057_ (.CLK(clknet_leaf_58_clk),
    .D(net1243),
    .RESET_B(_00102_),
    .Q(\mac_array.mac[11].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13058_ (.CLK(clknet_leaf_53_clk),
    .D(net2070),
    .RESET_B(_00103_),
    .Q(\mac_array.mac[11].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13059_ (.CLK(clknet_leaf_53_clk),
    .D(net2341),
    .RESET_B(_00104_),
    .Q(\mac_array.mac[11].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13060_ (.CLK(clknet_leaf_53_clk),
    .D(net2347),
    .RESET_B(_00105_),
    .Q(\mac_array.mac[11].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13061_ (.CLK(clknet_leaf_53_clk),
    .D(net2353),
    .RESET_B(_00106_),
    .Q(\mac_array.mac[11].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13062_ (.CLK(clknet_leaf_53_clk),
    .D(net2154),
    .RESET_B(_00107_),
    .Q(\mac_array.mac[11].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13063_ (.CLK(clknet_leaf_54_clk),
    .D(net2370),
    .RESET_B(_00108_),
    .Q(\mac_array.mac[11].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13064_ (.CLK(clknet_leaf_61_clk),
    .D(net2160),
    .RESET_B(_00109_),
    .Q(\mac_array.mac[10].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13065_ (.CLK(clknet_leaf_64_clk),
    .D(net1952),
    .RESET_B(_00110_),
    .Q(\mac_array.mac[10].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13066_ (.CLK(clknet_leaf_64_clk),
    .D(net1735),
    .RESET_B(_00111_),
    .Q(\mac_array.mac[10].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13067_ (.CLK(clknet_leaf_66_clk),
    .D(net2233),
    .RESET_B(_00112_),
    .Q(\mac_array.mac[10].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13068_ (.CLK(clknet_leaf_66_clk),
    .D(net1371),
    .RESET_B(_00113_),
    .Q(\mac_array.mac[10].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13069_ (.CLK(clknet_leaf_66_clk),
    .D(net2116),
    .RESET_B(_00114_),
    .Q(\mac_array.mac[10].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13070_ (.CLK(clknet_leaf_66_clk),
    .D(net2223),
    .RESET_B(_00115_),
    .Q(\mac_array.mac[10].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13071_ (.CLK(clknet_leaf_66_clk),
    .D(net1855),
    .RESET_B(_00116_),
    .Q(\mac_array.mac[10].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13072_ (.CLK(clknet_leaf_5_clk),
    .D(net1120),
    .RESET_B(_00117_),
    .Q(\mac_array.mac[9].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13073_ (.CLK(clknet_leaf_6_clk),
    .D(net1799),
    .RESET_B(_00118_),
    .Q(\mac_array.mac[9].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13074_ (.CLK(clknet_leaf_6_clk),
    .D(net1788),
    .RESET_B(_00119_),
    .Q(\mac_array.mac[9].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13075_ (.CLK(clknet_leaf_8_clk),
    .D(net1739),
    .RESET_B(_00120_),
    .Q(\mac_array.mac[9].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13076_ (.CLK(clknet_leaf_9_clk),
    .D(net1170),
    .RESET_B(_00121_),
    .Q(\mac_array.mac[9].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13077_ (.CLK(clknet_leaf_9_clk),
    .D(net1803),
    .RESET_B(_00122_),
    .Q(\mac_array.mac[9].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13078_ (.CLK(clknet_leaf_8_clk),
    .D(net1331),
    .RESET_B(_00123_),
    .Q(\mac_array.mac[9].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13079_ (.CLK(clknet_leaf_9_clk),
    .D(net1779),
    .RESET_B(_00124_),
    .Q(\mac_array.mac[9].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13080_ (.CLK(clknet_leaf_3_clk),
    .D(net1363),
    .RESET_B(_00125_),
    .Q(\mac_array.mac[8].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13081_ (.CLK(clknet_leaf_2_clk),
    .D(net2538),
    .RESET_B(_00126_),
    .Q(\mac_array.mac[8].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13082_ (.CLK(clknet_leaf_2_clk),
    .D(net2503),
    .RESET_B(_00127_),
    .Q(\mac_array.mac[8].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13083_ (.CLK(clknet_leaf_2_clk),
    .D(net2309),
    .RESET_B(_00128_),
    .Q(\mac_array.mac[8].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13084_ (.CLK(clknet_leaf_2_clk),
    .D(net1851),
    .RESET_B(_00129_),
    .Q(\mac_array.mac[8].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13085_ (.CLK(clknet_leaf_67_clk),
    .D(net1819),
    .RESET_B(_00130_),
    .Q(\mac_array.mac[8].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13086_ (.CLK(clknet_leaf_67_clk),
    .D(net1707),
    .RESET_B(_00131_),
    .Q(\mac_array.mac[8].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13087_ (.CLK(clknet_leaf_67_clk),
    .D(net1149),
    .RESET_B(_00132_),
    .Q(\mac_array.mac[8].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13088_ (.CLK(clknet_leaf_30_clk),
    .D(net2052),
    .RESET_B(_00133_),
    .Q(\mac_array.mac[7].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13089_ (.CLK(clknet_leaf_35_clk),
    .D(net2177),
    .RESET_B(_00134_),
    .Q(\mac_array.mac[7].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13090_ (.CLK(clknet_leaf_31_clk),
    .D(net1972),
    .RESET_B(_00135_),
    .Q(\mac_array.mac[7].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13091_ (.CLK(clknet_leaf_31_clk),
    .D(net2035),
    .RESET_B(_00136_),
    .Q(\mac_array.mac[7].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13092_ (.CLK(clknet_leaf_31_clk),
    .D(net1985),
    .RESET_B(_00137_),
    .Q(\mac_array.mac[7].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13093_ (.CLK(clknet_leaf_31_clk),
    .D(net1989),
    .RESET_B(_00138_),
    .Q(\mac_array.mac[7].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13094_ (.CLK(clknet_leaf_32_clk),
    .D(net1351),
    .RESET_B(_00139_),
    .Q(\mac_array.mac[7].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13095_ (.CLK(clknet_leaf_32_clk),
    .D(net2039),
    .RESET_B(_00140_),
    .Q(\mac_array.mac[7].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13096_ (.CLK(clknet_leaf_40_clk),
    .D(net2335),
    .RESET_B(_00141_),
    .Q(\mac_array.mac[6].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13097_ (.CLK(clknet_leaf_35_clk),
    .D(net1956),
    .RESET_B(_00142_),
    .Q(\mac_array.mac[6].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13098_ (.CLK(clknet_leaf_39_clk),
    .D(net2300),
    .RESET_B(_00143_),
    .Q(\mac_array.mac[6].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13099_ (.CLK(clknet_leaf_39_clk),
    .D(net2324),
    .RESET_B(_00144_),
    .Q(\mac_array.mac[6].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13100_ (.CLK(clknet_leaf_39_clk),
    .D(net2305),
    .RESET_B(_00145_),
    .Q(\mac_array.mac[6].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13101_ (.CLK(clknet_leaf_39_clk),
    .D(net1823),
    .RESET_B(_00146_),
    .Q(\mac_array.mac[6].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13102_ (.CLK(clknet_leaf_36_clk),
    .D(net2284),
    .RESET_B(_00147_),
    .Q(\mac_array.mac[6].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13103_ (.CLK(clknet_leaf_39_clk),
    .D(net2025),
    .RESET_B(_00148_),
    .Q(\mac_array.mac[6].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13104_ (.CLK(clknet_leaf_27_clk),
    .D(net2241),
    .RESET_B(_00149_),
    .Q(\mac_array.mac[5].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13105_ (.CLK(clknet_leaf_30_clk),
    .D(net2134),
    .RESET_B(_00150_),
    .Q(\mac_array.mac[5].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13106_ (.CLK(clknet_leaf_29_clk),
    .D(net2365),
    .RESET_B(_00151_),
    .Q(\mac_array.mac[5].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13107_ (.CLK(clknet_leaf_29_clk),
    .D(net1670),
    .RESET_B(_00152_),
    .Q(\mac_array.mac[5].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13108_ (.CLK(clknet_leaf_29_clk),
    .D(net2005),
    .RESET_B(_00153_),
    .Q(\mac_array.mac[5].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13109_ (.CLK(clknet_leaf_31_clk),
    .D(net2329),
    .RESET_B(_00154_),
    .Q(\mac_array.mac[5].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13110_ (.CLK(clknet_leaf_31_clk),
    .D(net1745),
    .RESET_B(_00155_),
    .Q(\mac_array.mac[5].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13111_ (.CLK(clknet_leaf_31_clk),
    .D(net1839),
    .RESET_B(_00156_),
    .Q(\mac_array.mac[5].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13112_ (.CLK(clknet_leaf_24_clk),
    .D(net2381),
    .RESET_B(_00157_),
    .Q(\mac_array.mac[4].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13113_ (.CLK(clknet_leaf_5_clk),
    .D(net1811),
    .RESET_B(_00158_),
    .Q(\mac_array.mac[4].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13114_ (.CLK(clknet_leaf_5_clk),
    .D(net2150),
    .RESET_B(_00159_),
    .Q(\mac_array.mac[4].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13115_ (.CLK(clknet_leaf_6_clk),
    .D(net2397),
    .RESET_B(_00160_),
    .Q(\mac_array.mac[4].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13116_ (.CLK(clknet_leaf_6_clk),
    .D(net2392),
    .RESET_B(_00161_),
    .Q(\mac_array.mac[4].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13117_ (.CLK(clknet_leaf_8_clk),
    .D(net1749),
    .RESET_B(_00162_),
    .Q(\mac_array.mac[4].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13118_ (.CLK(clknet_leaf_8_clk),
    .D(net2030),
    .RESET_B(_00163_),
    .Q(\mac_array.mac[4].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13119_ (.CLK(clknet_leaf_8_clk),
    .D(net1900),
    .RESET_B(_00164_),
    .Q(\mac_array.mac[4].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13120_ (.CLK(clknet_leaf_25_clk),
    .D(net2080),
    .RESET_B(_00165_),
    .Q(\mac_array.mac[3].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13121_ (.CLK(clknet_leaf_25_clk),
    .D(net1807),
    .RESET_B(_00166_),
    .Q(\mac_array.mac[3].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13122_ (.CLK(clknet_leaf_25_clk),
    .D(net2201),
    .RESET_B(_00167_),
    .Q(\mac_array.mac[3].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13123_ (.CLK(clknet_leaf_42_clk),
    .D(net2467),
    .RESET_B(_00168_),
    .Q(\mac_array.mac[3].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13124_ (.CLK(clknet_leaf_42_clk),
    .D(net2462),
    .RESET_B(_00169_),
    .Q(\mac_array.mac[3].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13125_ (.CLK(clknet_leaf_41_clk),
    .D(net1847),
    .RESET_B(_00170_),
    .Q(\mac_array.mac[3].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13126_ (.CLK(clknet_leaf_41_clk),
    .D(net2279),
    .RESET_B(_00171_),
    .Q(\mac_array.mac[3].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13127_ (.CLK(clknet_leaf_41_clk),
    .D(net1993),
    .RESET_B(_00172_),
    .Q(\mac_array.mac[3].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13128_ (.CLK(clknet_leaf_21_clk),
    .D(net1924),
    .RESET_B(_00173_),
    .Q(\mac_array.mac[2].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13129_ (.CLK(clknet_leaf_20_clk),
    .D(net1769),
    .RESET_B(_00174_),
    .Q(\mac_array.mac[2].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13130_ (.CLK(clknet_leaf_20_clk),
    .D(net1692),
    .RESET_B(_00175_),
    .Q(\mac_array.mac[2].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13131_ (.CLK(clknet_leaf_20_clk),
    .D(net2076),
    .RESET_B(_00176_),
    .Q(\mac_array.mac[2].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13132_ (.CLK(clknet_leaf_19_clk),
    .D(net1868),
    .RESET_B(_00177_),
    .Q(\mac_array.mac[2].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13133_ (.CLK(clknet_leaf_19_clk),
    .D(net1872),
    .RESET_B(_00178_),
    .Q(\mac_array.mac[2].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13134_ (.CLK(clknet_leaf_19_clk),
    .D(net1877),
    .RESET_B(_00179_),
    .Q(\mac_array.mac[2].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13135_ (.CLK(clknet_leaf_19_clk),
    .D(net1859),
    .RESET_B(_00180_),
    .Q(\mac_array.mac[2].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13136_ (.CLK(clknet_leaf_22_clk),
    .D(net1928),
    .RESET_B(_00181_),
    .Q(\mac_array.mac[1].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13137_ (.CLK(clknet_leaf_22_clk),
    .D(net1715),
    .RESET_B(_00182_),
    .Q(\mac_array.mac[1].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13138_ (.CLK(clknet_leaf_17_clk),
    .D(net1719),
    .RESET_B(_00183_),
    .Q(\mac_array.mac[1].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13139_ (.CLK(clknet_leaf_17_clk),
    .D(net2485),
    .RESET_B(_00184_),
    .Q(\mac_array.mac[1].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13140_ (.CLK(clknet_leaf_16_clk),
    .D(net2479),
    .RESET_B(_00185_),
    .Q(\mac_array.mac[1].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13141_ (.CLK(clknet_leaf_17_clk),
    .D(net1940),
    .RESET_B(_00186_),
    .Q(\mac_array.mac[1].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13142_ (.CLK(clknet_leaf_16_clk),
    .D(net2319),
    .RESET_B(_00187_),
    .Q(\mac_array.mac[1].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13143_ (.CLK(clknet_leaf_16_clk),
    .D(net1932),
    .RESET_B(_00188_),
    .Q(\mac_array.mac[1].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13144_ (.CLK(clknet_leaf_22_clk),
    .D(net2411),
    .RESET_B(_00189_),
    .Q(\mac_array.mac[0].mac_unit.b[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13145_ (.CLK(clknet_leaf_7_clk),
    .D(net2429),
    .RESET_B(_00190_),
    .Q(\mac_array.mac[0].mac_unit.b[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13146_ (.CLK(clknet_leaf_7_clk),
    .D(net2191),
    .RESET_B(_00191_),
    .Q(\mac_array.mac[0].mac_unit.b[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13147_ (.CLK(clknet_leaf_12_clk),
    .D(net2435),
    .RESET_B(_00192_),
    .Q(\mac_array.mac[0].mac_unit.b[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13148_ (.CLK(clknet_leaf_12_clk),
    .D(net2451),
    .RESET_B(_00193_),
    .Q(\mac_array.mac[0].mac_unit.b[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13149_ (.CLK(clknet_leaf_11_clk),
    .D(net1889),
    .RESET_B(_00194_),
    .Q(\mac_array.mac[0].mac_unit.b[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13150_ (.CLK(clknet_leaf_11_clk),
    .D(net1674),
    .RESET_B(_00195_),
    .Q(\mac_array.mac[0].mac_unit.b[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13151_ (.CLK(clknet_leaf_11_clk),
    .D(net1711),
    .RESET_B(_00196_),
    .Q(\mac_array.mac[0].mac_unit.b[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13152_ (.CLK(clknet_leaf_57_clk),
    .D(net1650),
    .RESET_B(_00197_),
    .Q(\line_buffer.data_out[120] ));
 sky130_fd_sc_hd__dfrtp_1 _13153_ (.CLK(clknet_leaf_57_clk),
    .D(net1335),
    .RESET_B(_00198_),
    .Q(\line_buffer.data_out[121] ));
 sky130_fd_sc_hd__dfrtp_1 _13154_ (.CLK(clknet_3_3__leaf_clk),
    .D(net1299),
    .RESET_B(_00199_),
    .Q(\line_buffer.data_out[122] ));
 sky130_fd_sc_hd__dfrtp_1 _13155_ (.CLK(clknet_leaf_57_clk),
    .D(net1367),
    .RESET_B(_00200_),
    .Q(\line_buffer.data_out[123] ));
 sky130_fd_sc_hd__dfrtp_1 _13156_ (.CLK(clknet_leaf_49_clk),
    .D(net2359),
    .RESET_B(_00201_),
    .Q(\line_buffer.data_out[124] ));
 sky130_fd_sc_hd__dfrtp_1 _13157_ (.CLK(clknet_leaf_49_clk),
    .D(net1124),
    .RESET_B(_00202_),
    .Q(\line_buffer.data_out[125] ));
 sky130_fd_sc_hd__dfrtp_1 _13158_ (.CLK(clknet_leaf_49_clk),
    .D(net1535),
    .RESET_B(_00203_),
    .Q(\line_buffer.data_out[126] ));
 sky130_fd_sc_hd__dfrtp_1 _13159_ (.CLK(clknet_leaf_49_clk),
    .D(net1454),
    .RESET_B(_00204_),
    .Q(\line_buffer.data_out[127] ));
 sky130_fd_sc_hd__dfrtp_1 _13160_ (.CLK(clknet_leaf_3_clk),
    .D(net1399),
    .RESET_B(_00205_),
    .Q(\result[11][0] ));
 sky130_fd_sc_hd__dfrtp_1 _13161_ (.CLK(clknet_leaf_3_clk),
    .D(net2574),
    .RESET_B(_00206_),
    .Q(\result[11][1] ));
 sky130_fd_sc_hd__dfrtp_1 _13162_ (.CLK(clknet_leaf_60_clk),
    .D(net1303),
    .RESET_B(_00207_),
    .Q(\result[11][2] ));
 sky130_fd_sc_hd__dfrtp_1 _13163_ (.CLK(clknet_leaf_60_clk),
    .D(net1319),
    .RESET_B(_00208_),
    .Q(\result[11][3] ));
 sky130_fd_sc_hd__dfrtp_1 _13164_ (.CLK(clknet_leaf_60_clk),
    .D(net2598),
    .RESET_B(_00209_),
    .Q(\result[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _13165_ (.CLK(clknet_leaf_60_clk),
    .D(net1327),
    .RESET_B(_00210_),
    .Q(\result[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _13166_ (.CLK(clknet_leaf_60_clk),
    .D(net1323),
    .RESET_B(_00211_),
    .Q(\result[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _13167_ (.CLK(clknet_leaf_4_clk),
    .D(net1235),
    .RESET_B(_00212_),
    .Q(\result[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _13168_ (.CLK(clknet_leaf_44_clk),
    .D(net1642),
    .RESET_B(_00213_),
    .Q(\line_buffer.data_out[112] ));
 sky130_fd_sc_hd__dfrtp_1 _13169_ (.CLK(clknet_leaf_44_clk),
    .D(net1831),
    .RESET_B(_00214_),
    .Q(\line_buffer.data_out[113] ));
 sky130_fd_sc_hd__dfrtp_1 _13170_ (.CLK(clknet_leaf_44_clk),
    .D(net2187),
    .RESET_B(_00215_),
    .Q(\line_buffer.data_out[114] ));
 sky130_fd_sc_hd__dfrtp_1 _13171_ (.CLK(clknet_leaf_46_clk),
    .D(net2403),
    .RESET_B(_00216_),
    .Q(\line_buffer.data_out[115] ));
 sky130_fd_sc_hd__dfrtp_1 _13172_ (.CLK(clknet_leaf_46_clk),
    .D(net2181),
    .RESET_B(_00217_),
    .Q(\line_buffer.data_out[116] ));
 sky130_fd_sc_hd__dfrtp_1 _13173_ (.CLK(clknet_leaf_47_clk),
    .D(net2211),
    .RESET_B(_00218_),
    .Q(\line_buffer.data_out[117] ));
 sky130_fd_sc_hd__dfrtp_1 _13174_ (.CLK(clknet_leaf_47_clk),
    .D(net1516),
    .RESET_B(_00219_),
    .Q(\line_buffer.data_out[118] ));
 sky130_fd_sc_hd__dfrtp_1 _13175_ (.CLK(clknet_leaf_47_clk),
    .D(net1502),
    .RESET_B(_00220_),
    .Q(\line_buffer.data_out[119] ));
 sky130_fd_sc_hd__dfrtp_1 _13176_ (.CLK(clknet_leaf_41_clk),
    .D(net1605),
    .RESET_B(_00221_),
    .Q(\line_buffer.data_out[104] ));
 sky130_fd_sc_hd__dfrtp_1 _13177_ (.CLK(clknet_leaf_42_clk),
    .D(net1759),
    .RESET_B(_00222_),
    .Q(\line_buffer.data_out[105] ));
 sky130_fd_sc_hd__dfrtp_1 _13178_ (.CLK(clknet_leaf_41_clk),
    .D(net1794),
    .RESET_B(_00223_),
    .Q(\line_buffer.data_out[106] ));
 sky130_fd_sc_hd__dfrtp_1 _13179_ (.CLK(clknet_leaf_42_clk),
    .D(net2260),
    .RESET_B(_00224_),
    .Q(\line_buffer.data_out[107] ));
 sky130_fd_sc_hd__dfrtp_1 _13180_ (.CLK(clknet_leaf_42_clk),
    .D(net2249),
    .RESET_B(_00225_),
    .Q(\line_buffer.data_out[108] ));
 sky130_fd_sc_hd__dfrtp_1 _13181_ (.CLK(clknet_leaf_41_clk),
    .D(net1162),
    .RESET_B(_00226_),
    .Q(\line_buffer.data_out[109] ));
 sky130_fd_sc_hd__dfrtp_1 _13182_ (.CLK(clknet_leaf_41_clk),
    .D(net1484),
    .RESET_B(_00227_),
    .Q(\line_buffer.data_out[110] ));
 sky130_fd_sc_hd__dfrtp_1 _13183_ (.CLK(clknet_leaf_41_clk),
    .D(net1387),
    .RESET_B(_00228_),
    .Q(\line_buffer.data_out[111] ));
 sky130_fd_sc_hd__dfrtp_1 _13184_ (.CLK(clknet_leaf_61_clk),
    .D(net1646),
    .RESET_B(_00229_),
    .Q(\line_buffer.data_out[96] ));
 sky130_fd_sc_hd__dfrtp_1 _13185_ (.CLK(clknet_leaf_61_clk),
    .D(net2058),
    .RESET_B(_00230_),
    .Q(\line_buffer.data_out[97] ));
 sky130_fd_sc_hd__dfrtp_1 _13186_ (.CLK(clknet_leaf_61_clk),
    .D(net2207),
    .RESET_B(_00231_),
    .Q(\line_buffer.data_out[98] ));
 sky130_fd_sc_hd__dfrtp_1 _13187_ (.CLK(clknet_leaf_61_clk),
    .D(net2592),
    .RESET_B(_00232_),
    .Q(\line_buffer.data_out[99] ));
 sky130_fd_sc_hd__dfrtp_1 _13188_ (.CLK(clknet_leaf_61_clk),
    .D(net2580),
    .RESET_B(_00233_),
    .Q(\line_buffer.data_out[100] ));
 sky130_fd_sc_hd__dfrtp_1 _13189_ (.CLK(clknet_leaf_61_clk),
    .D(net2586),
    .RESET_B(_00234_),
    .Q(\line_buffer.data_out[101] ));
 sky130_fd_sc_hd__dfrtp_1 _13190_ (.CLK(clknet_leaf_61_clk),
    .D(net1552),
    .RESET_B(_00235_),
    .Q(\line_buffer.data_out[102] ));
 sky130_fd_sc_hd__dfrtp_1 _13191_ (.CLK(clknet_leaf_61_clk),
    .D(net1498),
    .RESET_B(_00236_),
    .Q(\line_buffer.data_out[103] ));
 sky130_fd_sc_hd__dfrtp_1 _13192_ (.CLK(clknet_leaf_58_clk),
    .D(net1279),
    .RESET_B(_00237_),
    .Q(\line_buffer.data_out[88] ));
 sky130_fd_sc_hd__dfrtp_1 _13193_ (.CLK(clknet_leaf_58_clk),
    .D(net2140),
    .RESET_B(_00238_),
    .Q(\line_buffer.data_out[89] ));
 sky130_fd_sc_hd__dfrtp_1 _13194_ (.CLK(clknet_leaf_58_clk),
    .D(net2172),
    .RESET_B(_00239_),
    .Q(\line_buffer.data_out[90] ));
 sky130_fd_sc_hd__dfrtp_1 _13195_ (.CLK(clknet_leaf_58_clk),
    .D(net2295),
    .RESET_B(_00240_),
    .Q(\line_buffer.data_out[91] ));
 sky130_fd_sc_hd__dfrtp_1 _13196_ (.CLK(clknet_leaf_55_clk),
    .D(net2270),
    .RESET_B(_00241_),
    .Q(\line_buffer.data_out[92] ));
 sky130_fd_sc_hd__dfrtp_1 _13197_ (.CLK(clknet_leaf_55_clk),
    .D(net2289),
    .RESET_B(_00242_),
    .Q(\line_buffer.data_out[93] ));
 sky130_fd_sc_hd__dfrtp_1 _13198_ (.CLK(clknet_leaf_55_clk),
    .D(net1529),
    .RESET_B(_00243_),
    .Q(\line_buffer.data_out[94] ));
 sky130_fd_sc_hd__dfrtp_1 _13199_ (.CLK(clknet_leaf_55_clk),
    .D(net1458),
    .RESET_B(_00244_),
    .Q(\line_buffer.data_out[95] ));
 sky130_fd_sc_hd__dfrtp_1 _13200_ (.CLK(clknet_leaf_61_clk),
    .D(net1311),
    .RESET_B(_00245_),
    .Q(\line_buffer.data_out[80] ));
 sky130_fd_sc_hd__dfrtp_1 _13201_ (.CLK(clknet_leaf_0_clk),
    .D(net2064),
    .RESET_B(_00246_),
    .Q(\line_buffer.data_out[81] ));
 sky130_fd_sc_hd__dfrtp_1 _13202_ (.CLK(clknet_leaf_66_clk),
    .D(net2217),
    .RESET_B(_00247_),
    .Q(\line_buffer.data_out[82] ));
 sky130_fd_sc_hd__dfrtp_1 _13203_ (.CLK(clknet_leaf_66_clk),
    .D(net2112),
    .RESET_B(_00248_),
    .Q(\line_buffer.data_out[83] ));
 sky130_fd_sc_hd__dfrtp_1 _13204_ (.CLK(clknet_leaf_66_clk),
    .D(net2274),
    .RESET_B(_00249_),
    .Q(\line_buffer.data_out[84] ));
 sky130_fd_sc_hd__dfrtp_1 _13205_ (.CLK(clknet_leaf_66_clk),
    .D(net2473),
    .RESET_B(_00250_),
    .Q(\line_buffer.data_out[85] ));
 sky130_fd_sc_hd__dfrtp_1 _13206_ (.CLK(clknet_leaf_0_clk),
    .D(net1562),
    .RESET_B(_00251_),
    .Q(\line_buffer.data_out[86] ));
 sky130_fd_sc_hd__dfrtp_1 _13207_ (.CLK(clknet_leaf_66_clk),
    .D(net1506),
    .RESET_B(_00252_),
    .Q(\line_buffer.data_out[87] ));
 sky130_fd_sc_hd__dfrtp_1 _13208_ (.CLK(clknet_leaf_5_clk),
    .D(net1588),
    .RESET_B(_00253_),
    .Q(\line_buffer.data_out[72] ));
 sky130_fd_sc_hd__dfrtp_1 _13209_ (.CLK(clknet_leaf_8_clk),
    .D(net1660),
    .RESET_B(_00254_),
    .Q(\line_buffer.data_out[73] ));
 sky130_fd_sc_hd__dfrtp_1 _13210_ (.CLK(clknet_leaf_9_clk),
    .D(net1696),
    .RESET_B(_00255_),
    .Q(\line_buffer.data_out[74] ));
 sky130_fd_sc_hd__dfrtp_1 _13211_ (.CLK(clknet_leaf_9_clk),
    .D(net1976),
    .RESET_B(_00256_),
    .Q(\line_buffer.data_out[75] ));
 sky130_fd_sc_hd__dfrtp_1 _13212_ (.CLK(clknet_leaf_9_clk),
    .D(net2084),
    .RESET_B(_00257_),
    .Q(\line_buffer.data_out[76] ));
 sky130_fd_sc_hd__dfrtp_1 _13213_ (.CLK(clknet_leaf_9_clk),
    .D(net1885),
    .RESET_B(_00258_),
    .Q(\line_buffer.data_out[77] ));
 sky130_fd_sc_hd__dfrtp_1 _13214_ (.CLK(clknet_leaf_10_clk),
    .D(net1469),
    .RESET_B(_00259_),
    .Q(\line_buffer.data_out[78] ));
 sky130_fd_sc_hd__dfrtp_1 _13215_ (.CLK(clknet_leaf_10_clk),
    .D(net1413),
    .RESET_B(_00260_),
    .Q(\line_buffer.data_out[79] ));
 sky130_fd_sc_hd__dfrtp_1 _13216_ (.CLK(clknet_leaf_3_clk),
    .D(net1638),
    .RESET_B(_00261_),
    .Q(\line_buffer.data_out[64] ));
 sky130_fd_sc_hd__dfrtp_1 _13217_ (.CLK(clknet_leaf_1_clk),
    .D(net1948),
    .RESET_B(_00262_),
    .Q(\line_buffer.data_out[65] ));
 sky130_fd_sc_hd__dfrtp_1 _13218_ (.CLK(clknet_leaf_1_clk),
    .D(net1962),
    .RESET_B(_00263_),
    .Q(\line_buffer.data_out[66] ));
 sky130_fd_sc_hd__dfrtp_1 _13219_ (.CLK(clknet_leaf_1_clk),
    .D(net2313),
    .RESET_B(_00264_),
    .Q(\line_buffer.data_out[67] ));
 sky130_fd_sc_hd__dfrtp_1 _13220_ (.CLK(clknet_leaf_1_clk),
    .D(net1666),
    .RESET_B(_00265_),
    .Q(\line_buffer.data_out[68] ));
 sky130_fd_sc_hd__dfrtp_1 _13221_ (.CLK(clknet_leaf_1_clk),
    .D(net1765),
    .RESET_B(_00266_),
    .Q(\line_buffer.data_out[69] ));
 sky130_fd_sc_hd__dfrtp_1 _13222_ (.CLK(clknet_leaf_1_clk),
    .D(net1543),
    .RESET_B(_00267_),
    .Q(\line_buffer.data_out[70] ));
 sky130_fd_sc_hd__dfrtp_1 _13223_ (.CLK(clknet_leaf_1_clk),
    .D(net1494),
    .RESET_B(_00268_),
    .Q(\line_buffer.data_out[71] ));
 sky130_fd_sc_hd__dfrtp_1 _13224_ (.CLK(clknet_leaf_30_clk),
    .D(net1617),
    .RESET_B(_00269_),
    .Q(\line_buffer.data_out[56] ));
 sky130_fd_sc_hd__dfrtp_1 _13225_ (.CLK(clknet_leaf_30_clk),
    .D(net1936),
    .RESET_B(_00270_),
    .Q(\line_buffer.data_out[57] ));
 sky130_fd_sc_hd__dfrtp_1 _13226_ (.CLK(clknet_leaf_30_clk),
    .D(net1911),
    .RESET_B(_00271_),
    .Q(\line_buffer.data_out[58] ));
 sky130_fd_sc_hd__dfrtp_1 _13227_ (.CLK(clknet_leaf_34_clk),
    .D(net1359),
    .RESET_B(_00272_),
    .Q(\line_buffer.data_out[59] ));
 sky130_fd_sc_hd__dfrtp_1 _13228_ (.CLK(clknet_leaf_34_clk),
    .D(net2254),
    .RESET_B(_00273_),
    .Q(\line_buffer.data_out[60] ));
 sky130_fd_sc_hd__dfrtp_1 _13229_ (.CLK(clknet_leaf_34_clk),
    .D(net2375),
    .RESET_B(_00274_),
    .Q(\line_buffer.data_out[61] ));
 sky130_fd_sc_hd__dfrtp_1 _13230_ (.CLK(clknet_leaf_34_clk),
    .D(net1478),
    .RESET_B(_00275_),
    .Q(\line_buffer.data_out[62] ));
 sky130_fd_sc_hd__dfrtp_1 _13231_ (.CLK(clknet_leaf_34_clk),
    .D(net1440),
    .RESET_B(_00276_),
    .Q(\line_buffer.data_out[63] ));
 sky130_fd_sc_hd__dfrtp_1 _13232_ (.CLK(clknet_leaf_27_clk),
    .D(net1628),
    .RESET_B(_00277_),
    .Q(\line_buffer.data_out[48] ));
 sky130_fd_sc_hd__dfrtp_1 _13233_ (.CLK(clknet_leaf_27_clk),
    .D(net1981),
    .RESET_B(_00278_),
    .Q(\line_buffer.data_out[49] ));
 sky130_fd_sc_hd__dfrtp_1 _13234_ (.CLK(clknet_leaf_40_clk),
    .D(net2021),
    .RESET_B(_00279_),
    .Q(\line_buffer.data_out[50] ));
 sky130_fd_sc_hd__dfrtp_1 _13235_ (.CLK(clknet_leaf_36_clk),
    .D(net2445),
    .RESET_B(_00280_),
    .Q(\line_buffer.data_out[51] ));
 sky130_fd_sc_hd__dfrtp_1 _13236_ (.CLK(clknet_leaf_36_clk),
    .D(net2440),
    .RESET_B(_00281_),
    .Q(\line_buffer.data_out[52] ));
 sky130_fd_sc_hd__dfrtp_1 _13237_ (.CLK(clknet_leaf_36_clk),
    .D(net2237),
    .RESET_B(_00282_),
    .Q(\line_buffer.data_out[53] ));
 sky130_fd_sc_hd__dfrtp_1 _13238_ (.CLK(clknet_leaf_36_clk),
    .D(net1512),
    .RESET_B(_00283_),
    .Q(\line_buffer.data_out[54] ));
 sky130_fd_sc_hd__dfrtp_1 _13239_ (.CLK(clknet_leaf_36_clk),
    .D(net1409),
    .RESET_B(_00284_),
    .Q(\line_buffer.data_out[55] ));
 sky130_fd_sc_hd__dfrtp_1 _13240_ (.CLK(clknet_leaf_30_clk),
    .D(net1613),
    .RESET_B(_00285_),
    .Q(\line_buffer.data_out[40] ));
 sky130_fd_sc_hd__dfrtp_1 _13241_ (.CLK(clknet_leaf_30_clk),
    .D(net1723),
    .RESET_B(_00286_),
    .Q(\line_buffer.data_out[41] ));
 sky130_fd_sc_hd__dfrtp_1 _13242_ (.CLK(clknet_leaf_31_clk),
    .D(net1815),
    .RESET_B(_00287_),
    .Q(\line_buffer.data_out[42] ));
 sky130_fd_sc_hd__dfrtp_1 _13243_ (.CLK(clknet_leaf_31_clk),
    .D(net2245),
    .RESET_B(_00288_),
    .Q(\line_buffer.data_out[43] ));
 sky130_fd_sc_hd__dfrtp_1 _13244_ (.CLK(clknet_leaf_29_clk),
    .D(net1997),
    .RESET_B(_00289_),
    .Q(\line_buffer.data_out[44] ));
 sky130_fd_sc_hd__dfrtp_1 _13245_ (.CLK(clknet_leaf_29_clk),
    .D(net1158),
    .RESET_B(_00290_),
    .Q(\line_buffer.data_out[45] ));
 sky130_fd_sc_hd__dfrtp_1 _13246_ (.CLK(clknet_leaf_29_clk),
    .D(net1473),
    .RESET_B(_00291_),
    .Q(\line_buffer.data_out[46] ));
 sky130_fd_sc_hd__dfrtp_1 _13247_ (.CLK(clknet_leaf_31_clk),
    .D(net1423),
    .RESET_B(_00292_),
    .Q(\line_buffer.data_out[47] ));
 sky130_fd_sc_hd__dfrtp_1 _13248_ (.CLK(clknet_leaf_5_clk),
    .D(net1592),
    .RESET_B(_00293_),
    .Q(\line_buffer.data_out[32] ));
 sky130_fd_sc_hd__dfrtp_1 _13249_ (.CLK(clknet_leaf_6_clk),
    .D(net1679),
    .RESET_B(_00294_),
    .Q(\line_buffer.data_out[33] ));
 sky130_fd_sc_hd__dfrtp_1 _13250_ (.CLK(clknet_leaf_6_clk),
    .D(net1701),
    .RESET_B(_00295_),
    .Q(\line_buffer.data_out[34] ));
 sky130_fd_sc_hd__dfrtp_1 _13251_ (.CLK(clknet_leaf_6_clk),
    .D(net2520),
    .RESET_B(_00296_),
    .Q(\line_buffer.data_out[35] ));
 sky130_fd_sc_hd__dfrtp_1 _13252_ (.CLK(clknet_leaf_8_clk),
    .D(net2227),
    .RESET_B(_00297_),
    .Q(\line_buffer.data_out[36] ));
 sky130_fd_sc_hd__dfrtp_1 _13253_ (.CLK(clknet_leaf_8_clk),
    .D(net2515),
    .RESET_B(_00298_),
    .Q(\line_buffer.data_out[37] ));
 sky130_fd_sc_hd__dfrtp_1 _13254_ (.CLK(clknet_leaf_8_clk),
    .D(net1405),
    .RESET_B(_00299_),
    .Q(\line_buffer.data_out[38] ));
 sky130_fd_sc_hd__dfrtp_1 _13255_ (.CLK(clknet_leaf_8_clk),
    .D(net1383),
    .RESET_B(_00300_),
    .Q(\line_buffer.data_out[39] ));
 sky130_fd_sc_hd__dfrtp_1 _13256_ (.CLK(clknet_leaf_42_clk),
    .D(net1609),
    .RESET_B(_00301_),
    .Q(\line_buffer.data_out[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13257_ (.CLK(clknet_leaf_42_clk),
    .D(net1754),
    .RESET_B(_00302_),
    .Q(\line_buffer.data_out[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13258_ (.CLK(clknet_leaf_41_clk),
    .D(net1784),
    .RESET_B(_00303_),
    .Q(\line_buffer.data_out[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13259_ (.CLK(clknet_leaf_38_clk),
    .D(net1174),
    .RESET_B(_00304_),
    .Q(\line_buffer.data_out[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13260_ (.CLK(clknet_leaf_38_clk),
    .D(net1096),
    .RESET_B(_00305_),
    .Q(\line_buffer.data_out[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13261_ (.CLK(clknet_leaf_38_clk),
    .D(net2423),
    .RESET_B(_00306_),
    .Q(\line_buffer.data_out[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13262_ (.CLK(clknet_leaf_38_clk),
    .D(net1347),
    .RESET_B(_00307_),
    .Q(\line_buffer.data_out[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13263_ (.CLK(clknet_leaf_38_clk),
    .D(net1427),
    .RESET_B(_00308_),
    .Q(\line_buffer.data_out[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13264_ (.CLK(clknet_leaf_20_clk),
    .D(net1634),
    .RESET_B(_00309_),
    .Q(\line_buffer.data_out[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13265_ (.CLK(clknet_leaf_19_clk),
    .D(net1775),
    .RESET_B(_00310_),
    .Q(\line_buffer.data_out[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13266_ (.CLK(clknet_leaf_18_clk),
    .D(net1968),
    .RESET_B(_00311_),
    .Q(\line_buffer.data_out[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13267_ (.CLK(clknet_leaf_19_clk),
    .D(net1881),
    .RESET_B(_00312_),
    .Q(\line_buffer.data_out[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13268_ (.CLK(clknet_leaf_19_clk),
    .D(net2264),
    .RESET_B(_00313_),
    .Q(\line_buffer.data_out[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13269_ (.CLK(clknet_leaf_19_clk),
    .D(net2387),
    .RESET_B(_00314_),
    .Q(\line_buffer.data_out[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13270_ (.CLK(clknet_leaf_19_clk),
    .D(net1436),
    .RESET_B(_00315_),
    .Q(\line_buffer.data_out[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13271_ (.CLK(clknet_leaf_19_clk),
    .D(net1395),
    .RESET_B(_00316_),
    .Q(\line_buffer.data_out[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13272_ (.CLK(clknet_leaf_22_clk),
    .D(net1572),
    .RESET_B(_00317_),
    .Q(\line_buffer.data_out[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13273_ (.CLK(clknet_leaf_17_clk),
    .D(net1906),
    .RESET_B(_00318_),
    .Q(\line_buffer.data_out[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13274_ (.CLK(clknet_leaf_17_clk),
    .D(net1283),
    .RESET_B(_00319_),
    .Q(\line_buffer.data_out[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13275_ (.CLK(clknet_leaf_16_clk),
    .D(net1827),
    .RESET_B(_00320_),
    .Q(\line_buffer.data_out[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13276_ (.CLK(clknet_leaf_16_clk),
    .D(net2103),
    .RESET_B(_00321_),
    .Q(\line_buffer.data_out[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13277_ (.CLK(clknet_leaf_16_clk),
    .D(net2457),
    .RESET_B(_00322_),
    .Q(\line_buffer.data_out[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13278_ (.CLK(clknet_leaf_18_clk),
    .D(net1463),
    .RESET_B(_00323_),
    .Q(\line_buffer.data_out[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13279_ (.CLK(clknet_leaf_18_clk),
    .D(net1431),
    .RESET_B(_00324_),
    .Q(\line_buffer.data_out[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13280_ (.CLK(clknet_leaf_22_clk),
    .D(net1576),
    .RESET_B(_00325_),
    .Q(\line_buffer.data_out[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13281_ (.CLK(clknet_leaf_11_clk),
    .D(net1654),
    .RESET_B(_00326_),
    .Q(\line_buffer.data_out[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13282_ (.CLK(clknet_leaf_11_clk),
    .D(net1688),
    .RESET_B(_00327_),
    .Q(\line_buffer.data_out[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13283_ (.CLK(clknet_leaf_11_clk),
    .D(net1863),
    .RESET_B(_00328_),
    .Q(\line_buffer.data_out[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13284_ (.CLK(clknet_leaf_13_clk),
    .D(net2491),
    .RESET_B(_00329_),
    .Q(\line_buffer.data_out[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13285_ (.CLK(clknet_leaf_13_clk),
    .D(net2497),
    .RESET_B(_00330_),
    .Q(\line_buffer.data_out[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13286_ (.CLK(clknet_leaf_13_clk),
    .D(net1490),
    .RESET_B(_00331_),
    .Q(\line_buffer.data_out[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13287_ (.CLK(clknet_leaf_13_clk),
    .D(net1450),
    .RESET_B(_00332_),
    .Q(\line_buffer.data_out[7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 fanout100 (.A(net1531),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 fanout101 (.A(net2656),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 fanout102 (.A(net2355),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net1365),
    .X(net103));
 sky130_fd_sc_hd__buf_4 fanout104 (.A(net1297),
    .X(net104));
 sky130_fd_sc_hd__buf_4 fanout105 (.A(net1333),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 fanout106 (.A(net2447),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 fanout107 (.A(net2431),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 fanout108 (.A(net2425),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 fanout109 (.A(net2007),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 fanout110 (.A(net2315),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 fanout111 (.A(net2475),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 fanout112 (.A(net2481),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 fanout113 (.A(net2798),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 fanout114 (.A(net2869),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 fanout115 (.A(net2072),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 fanout116 (.A(net2808),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 fanout117 (.A(net2276),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 fanout118 (.A(net2459),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 fanout119 (.A(net2464),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 fanout120 (.A(net2027),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 fanout121 (.A(net2389),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 fanout122 (.A(net2394),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 fanout123 (.A(net2377),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 fanout124 (.A(net1741),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 fanout125 (.A(net2838),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 fanout126 (.A(net2361),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 fanout127 (.A(net2281),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 fanout128 (.A(net781),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 fanout129 (.A(net1003),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 fanout130 (.A(net2297),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 fanout131 (.A(net2331),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net1349),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 fanout133 (.A(net991),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 fanout134 (.A(net1006),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 fanout135 (.A(net1009),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 fanout136 (.A(net1703),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 fanout137 (.A(net2499),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 fanout138 (.A(net2534),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net1361),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net1329),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 fanout141 (.A(net2824),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 fanout142 (.A(net2773),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 fanout143 (.A(net2819),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 fanout144 (.A(net2219),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net1369),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 fanout146 (.A(net2229),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 fanout147 (.A(net2156),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 fanout148 (.A(net2768),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 fanout149 (.A(net2349),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 fanout150 (.A(net2343),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 fanout151 (.A(net2337),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 fanout152 (.A(net2066),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net1241),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 fanout154 (.A(net2505),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 fanout155 (.A(net2413),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 fanout156 (.A(net2522),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 fanout157 (.A(net2528),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 fanout158 (.A(net2540),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 fanout159 (.A(net2803),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 fanout160 (.A(net3010),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 fanout161 (.A(net2970),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 fanout162 (.A(net2142),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net1353),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 fanout164 (.A(net2852),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 fanout165 (.A(net2105),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(net2367),
    .X(net166));
 sky130_fd_sc_hd__buf_6 fanout167 (.A(net1874),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(net2326),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(net1681),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(net2032),
    .X(net170));
 sky130_fd_sc_hd__buf_6 fanout171 (.A(net2086),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net1796),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net1921),
    .X(net173));
 sky130_fd_sc_hd__buf_12 fanout174 (.A(net1377),
    .X(net174));
 sky130_fd_sc_hd__buf_12 fanout175 (.A(net1389),
    .X(net175));
 sky130_fd_sc_hd__buf_6 fanout176 (.A(net2286),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(net2606),
    .X(net177));
 sky130_fd_sc_hd__buf_6 fanout178 (.A(net2611),
    .X(net178));
 sky130_fd_sc_hd__buf_12 fanout179 (.A(net1554),
    .X(net179));
 sky130_fd_sc_hd__buf_12 fanout180 (.A(net1564),
    .X(net180));
 sky130_fd_sc_hd__buf_8 fanout181 (.A(net1373),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 fanout182 (.A(net2162),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 fanout183 (.A(net2127),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 fanout184 (.A(net2118),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 fanout185 (.A(net2193),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 fanout186 (.A(net2095),
    .X(net186));
 sky130_fd_sc_hd__buf_8 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_8 fanout188 (.A(net195),
    .X(net188));
 sky130_fd_sc_hd__buf_8 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_8 fanout190 (.A(net195),
    .X(net190));
 sky130_fd_sc_hd__buf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_8 fanout192 (.A(net195),
    .X(net192));
 sky130_fd_sc_hd__buf_8 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_8 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_12 fanout195 (.A(net1),
    .X(net195));
 sky130_fd_sc_hd__buf_8 fanout196 (.A(net210),
    .X(net196));
 sky130_fd_sc_hd__buf_8 fanout197 (.A(net210),
    .X(net197));
 sky130_fd_sc_hd__buf_8 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_8 fanout199 (.A(net210),
    .X(net199));
 sky130_fd_sc_hd__buf_8 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_8 fanout201 (.A(net210),
    .X(net201));
 sky130_fd_sc_hd__buf_8 fanout202 (.A(net210),
    .X(net202));
 sky130_fd_sc_hd__buf_8 fanout203 (.A(net206),
    .X(net203));
 sky130_fd_sc_hd__buf_6 fanout204 (.A(net206),
    .X(net204));
 sky130_fd_sc_hd__buf_8 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_8 fanout206 (.A(net210),
    .X(net206));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_8 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_8 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_8 fanout210 (.A(net1),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(net1247),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout35 (.A(net1247),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(net1246),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(net250),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 fanout38 (.A(net1486),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 fanout39 (.A(net2493),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 fanout40 (.A(net2487),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 fanout41 (.A(net2792),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 fanout42 (.A(net2453),
    .X(net42));
 sky130_fd_sc_hd__buf_4 fanout43 (.A(net1281),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 fanout44 (.A(net1902),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 fanout45 (.A(net1568),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 fanout46 (.A(net2813),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 fanout47 (.A(net2383),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 fanout48 (.A(net1964),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 fanout49 (.A(net1771),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 fanout50 (.A(net1630),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net1345),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 fanout52 (.A(net2419),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 fanout53 (.A(net2846),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 fanout54 (.A(net1781),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 fanout55 (.A(net1751),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 fanout56 (.A(net2950),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 fanout57 (.A(net2511),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 fanout58 (.A(net2517),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 fanout59 (.A(net1698),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 fanout60 (.A(net1676),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 fanout61 (.A(net1508),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 fanout62 (.A(net3346),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 fanout63 (.A(net2442),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 fanout64 (.A(net964),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 fanout65 (.A(net967),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 fanout66 (.A(net556),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 fanout67 (.A(net796),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 fanout68 (.A(net2251),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(net1357),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 fanout70 (.A(net916),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 fanout71 (.A(net1761),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 fanout72 (.A(net1662),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 fanout73 (.A(net1958),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 fanout74 (.A(net1465),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 fanout75 (.A(net1656),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 fanout76 (.A(net1584),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 fanout77 (.A(net1558),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 fanout78 (.A(net2469),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 fanout79 (.A(net2213),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 fanout80 (.A(net2060),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(net1309),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 fanout82 (.A(net1525),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 fanout83 (.A(net2829),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 fanout84 (.A(net2266),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 fanout85 (.A(net2291),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 fanout86 (.A(net2168),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 fanout87 (.A(net2136),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(net1277),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 fanout89 (.A(net2582),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 fanout90 (.A(net2576),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 fanout91 (.A(net2588),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 fanout92 (.A(net2203),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 fanout93 (.A(net2054),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 fanout94 (.A(net1480),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 fanout95 (.A(net2256),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 fanout96 (.A(net1790),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 fanout97 (.A(net1756),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 fanout98 (.A(net2399),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 fanout99 (.A(net2183),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net2726),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net2748),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net1302),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(net2879),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(net2881),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(net2882),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(net262),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(net3250),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(net1078),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(net237),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(net1079),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_00355_),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(net256),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net2989),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(net2884),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(net2886),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(net2887),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(net258),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(net2889),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(net2891),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(net2892),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(net260),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(net2903),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(net2905),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net1314),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_00381_),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(net264),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(net2911),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(net2913),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_00544_),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(net268),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(net2906),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(net2908),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(net2909),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(net266),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net2993),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(net2898),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(net2900),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(net2901),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(net270),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(net3129),
    .X(net1244));
 sky130_fd_sc_hd__clkbuf_4 hold1035 (.A(net249),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_00693_),
    .X(net1246));
 sky130_fd_sc_hd__clkbuf_4 hold1037 (.A(net36),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(net2897),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(net272),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net1294),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(net2914),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(net2916),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(net2917),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(net280),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(net2919),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(net2921),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(net2922),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(net278),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(net2924),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(net2926),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net2985),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(net2927),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(net274),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\result[0][7] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(net1137),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(net281),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(net1138),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_00365_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(net282),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(net2928),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(net2930),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net1318),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(net2931),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(net284),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(net2955),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(net2957),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_00380_),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(net288),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(net2940),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(net289),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(net2944),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(net290),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net3016),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(net2958),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(net285),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(net2962),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(net286),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(net2932),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(net2934),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(net2935),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(net292),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(net2946),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(net2948),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net1322),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_00373_),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(net294),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(net2992),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(net2994),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_00379_),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(net314),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(net2975),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(net303),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(net2978),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(net304),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net3019),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(net2980),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(net2982),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(net2983),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(net310),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(net3005),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(net3007),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(net3008),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(net306),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(net2999),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(net307),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net1046),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net1326),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(net3003),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(net308),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(net2988),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(net2990),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(net2991),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(net312),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(net2984),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(net2986),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(net2987),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(net316),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net3035),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(net3015),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(net3017),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_00543_),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(net318),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(net3018),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(net3020),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_00542_),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(net320),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(net3034),
    .X(net1328));
 sky130_fd_sc_hd__buf_1 hold1119 (.A(net321),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net3039),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(net3038),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(net322),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(net3028),
    .X(net1332));
 sky130_fd_sc_hd__buf_1 hold1123 (.A(net323),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(net3032),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(net324),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(net3025),
    .X(net1336));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1127 (.A(net3027),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_00406_),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(net328),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net1332),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(net2784),
    .X(net1340));
 sky130_fd_sc_hd__clkbuf_2 hold1131 (.A(net2786),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_00397_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(net326),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(net3040),
    .X(net1344));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1135 (.A(net338),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(net3044),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(net3046),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\mac_array.mac[7].mac_unit.b[6] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(net340),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net3033),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(net3051),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(net341),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(net3053),
    .X(net1352));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1143 (.A(net357),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(net3057),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(net358),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(net3059),
    .X(net1356));
 sky130_fd_sc_hd__buf_1 hold1147 (.A(net352),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(net3061),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(net353),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net2785),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(net3063),
    .X(net1360));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1151 (.A(net3065),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(net3066),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(net368),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(net3073),
    .X(net1364));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1155 (.A(net369),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_00532_),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(net370),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(net3067),
    .X(net1368));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1159 (.A(net374),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net1342),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(net3071),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(net375),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(net3081),
    .X(net1372));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1163 (.A(net3083),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_00386_),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(net381),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(net3084),
    .X(net1376));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1167 (.A(net3086),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_00393_),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(net395),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net3026),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(net3089),
    .X(net1380));
 sky130_fd_sc_hd__buf_4 hold1171 (.A(net405),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_00632_),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(net406),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(net3599),
    .X(net1384));
 sky130_fd_sc_hd__buf_4 hold1175 (.A(net412),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(net3087),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(net413),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(net3091),
    .X(net1388));
 sky130_fd_sc_hd__buf_1 hold1179 (.A(net3093),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net1338),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_00392_),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(net404),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(net3094),
    .X(net1392));
 sky130_fd_sc_hd__buf_4 hold1183 (.A(net414),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(net3096),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(net415),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(net3660),
    .X(net1396));
 sky130_fd_sc_hd__clkbuf_2 hold1187 (.A(net333),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(net2783),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(net334),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net3622),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(net1441),
    .X(net1400));
 sky130_fd_sc_hd__buf_1 hold1191 (.A(net1443),
    .X(net1401));
 sky130_fd_sc_hd__clkbuf_2 hold1192 (.A(_00670_),
    .X(net1402));
 sky130_fd_sc_hd__clkbuf_4 hold1193 (.A(_00679_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(net2952),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(net2954),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(net3105),
    .X(net1406));
 sky130_fd_sc_hd__buf_4 hold1197 (.A(net423),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(net3107),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(net424),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net2751),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net2680),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(net3117),
    .X(net1410));
 sky130_fd_sc_hd__clkbuf_4 hold1201 (.A(net427),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(net3119),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(net428),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\result[13][3] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(net344),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_06100_),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(net345),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(net3191),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(net346),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net3399),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(net3109),
    .X(net1420));
 sky130_fd_sc_hd__buf_4 hold1211 (.A(net429),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(net3111),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(net430),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(net3113),
    .X(net1424));
 sky130_fd_sc_hd__buf_4 hold1215 (.A(net433),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(net3115),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(net434),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(net3121),
    .X(net1428));
 sky130_fd_sc_hd__clkbuf_4 hold1219 (.A(net437),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(net2822),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_00656_),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(net438),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(net1618),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(net1620),
    .X(net1433));
 sky130_fd_sc_hd__clkbuf_4 hold1224 (.A(_00675_),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(net2815),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(net2817),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(net3123),
    .X(net1437));
 sky130_fd_sc_hd__buf_4 hold1228 (.A(net442),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(net3127),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net3661),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(net443),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\control_fsm.line_write_addr[0] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(net1400),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(net342),
    .X(net1443));
 sky130_fd_sc_hd__clkbuf_2 hold1234 (.A(net1401),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(_00382_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(net343),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(net3141),
    .X(net1447));
 sky130_fd_sc_hd__buf_4 hold1238 (.A(net452),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(net3143),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net1398),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(net453),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(net3131),
    .X(net1451));
 sky130_fd_sc_hd__buf_4 hold1242 (.A(net457),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(_00536_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(net458),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(net3133),
    .X(net1455));
 sky130_fd_sc_hd__buf_4 hold1246 (.A(net470),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(net3135),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(net471),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(net3145),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net2843),
    .X(net335));
 sky130_fd_sc_hd__buf_2 hold1250 (.A(net3147),
    .X(net1460));
 sky130_fd_sc_hd__clkbuf_4 hold1251 (.A(_00673_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(net2794),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(net2796),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(net3567),
    .X(net1464));
 sky130_fd_sc_hd__buf_1 hold1255 (.A(net481),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(net74),
    .X(net1466));
 sky130_fd_sc_hd__buf_1 hold1257 (.A(net3579),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_00591_),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(net483),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_03270_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(net3137),
    .X(net1470));
 sky130_fd_sc_hd__buf_4 hold1261 (.A(net508),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(net3139),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(net509),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(net3788),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\line_buffer.data_out[34] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(net3153),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(net558),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\line_buffer.data_out[110] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net1547),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(net536),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(net94),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(net537),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(_00559_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(net538),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(net3746),
    .X(net1485));
 sky130_fd_sc_hd__buf_1 hold1276 (.A(net539),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(net38),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(net540),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(_00663_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net3041),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(net541),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(net3160),
    .X(net1491));
 sky130_fd_sc_hd__buf_4 hold1282 (.A(net550),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(_00600_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(net551),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(net3164),
    .X(net1495));
 sky130_fd_sc_hd__clkbuf_4 hold1286 (.A(net534),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(_00568_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(net535),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(net3154),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net3045),
    .X(net339));
 sky130_fd_sc_hd__buf_4 hold1290 (.A(net597),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(_00552_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(net598),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(net3162),
    .X(net1503));
 sky130_fd_sc_hd__buf_4 hold1294 (.A(net622),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(_00584_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(net623),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\line_buffer.data_out[54] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(net613),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(net61),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net2763),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net1348),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(net614),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(_00615_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(net615),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(net3166),
    .X(net1513));
 sky130_fd_sc_hd__clkbuf_4 hold1304 (.A(net490),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(_00551_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(net491),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(net3363),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(net1191),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(net388),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net3052),
    .X(net341));
 sky130_fd_sc_hd__buf_1 hold1310 (.A(net1192),
    .X(net1520));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1311 (.A(net3367),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_00384_),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(net366),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(net3827),
    .X(net1524));
 sky130_fd_sc_hd__buf_1 hold1315 (.A(net696),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(net82),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(net697),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_00575_),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(net698),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net1442),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(net3826),
    .X(net1530));
 sky130_fd_sc_hd__clkbuf_2 hold1321 (.A(net701),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(net100),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(net702),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_00535_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(net703),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(net2863),
    .X(net1536));
 sky130_fd_sc_hd__buf_2 hold1327 (.A(net2865),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_00407_),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(net379),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net1445),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(net3195),
    .X(net1540));
 sky130_fd_sc_hd__buf_4 hold1331 (.A(net628),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_00599_),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(net629),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(net2842),
    .X(net1544));
 sky130_fd_sc_hd__clkbuf_2 hold1335 (.A(net2844),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_03269_),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(_00396_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(net337),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(net3197),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net1414),
    .X(net344));
 sky130_fd_sc_hd__buf_4 hold1340 (.A(net650),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(_00567_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(net651),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(net3199),
    .X(net1553));
 sky130_fd_sc_hd__clkbuf_2 hold1344 (.A(net3201),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(_00388_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(net399),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\line_buffer.data_out[86] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(net724),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(net77),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net1416),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(net725),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(_00583_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(net726),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(net3202),
    .X(net1563));
 sky130_fd_sc_hd__clkbuf_2 hold1354 (.A(net3204),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(_00387_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(net411),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\line_buffer.data_out[8] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(net730),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(net3794),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net1418),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(_00649_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(net732),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(net3206),
    .X(net1573));
 sky130_fd_sc_hd__buf_4 hold1364 (.A(net677),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(_00657_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(net678),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\control_fsm.state[2] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(net359),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(net246),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net2545),
    .X(net347));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1370 (.A(net360),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(_00408_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(net361),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\line_buffer.data_out[72] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(net760),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(net76),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(net761),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(_00585_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(net762),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(net3223),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net2547),
    .X(net348));
 sky130_fd_sc_hd__buf_4 hold1380 (.A(net502),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(_00625_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(net503),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\control_fsm.state[0] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(net1197),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(net254),
    .X(net1595));
 sky130_fd_sc_hd__buf_1 hold1386 (.A(net1198),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(_03266_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(net2404),
    .X(net1598));
 sky130_fd_sc_hd__clkbuf_2 hold1389 (.A(net2406),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net2549),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_00395_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(net419),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(net3231),
    .X(net1602));
 sky130_fd_sc_hd__buf_4 hold1393 (.A(net605),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(_00553_),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(net606),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(net3227),
    .X(net1606));
 sky130_fd_sc_hd__buf_4 hold1397 (.A(net644),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_00633_),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(net645),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net1070),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net3473),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(net3233),
    .X(net1610));
 sky130_fd_sc_hd__clkbuf_4 hold1401 (.A(net494),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(_00617_),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(net495),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(net3663),
    .X(net1614));
 sky130_fd_sc_hd__clkbuf_4 hold1405 (.A(net520),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(net3239),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(net521),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\control_fsm.line_write_addr[3] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(net1432),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net2974),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(net400),
    .X(net1620));
 sky130_fd_sc_hd__clkbuf_2 hold1411 (.A(net1433),
    .X(net1621));
 sky130_fd_sc_hd__buf_4 hold1412 (.A(_00688_),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(_00385_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(net402),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(net3240),
    .X(net1625));
 sky130_fd_sc_hd__buf_4 hold1416 (.A(net530),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(_00609_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(net531),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\line_buffer.data_out[16] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net1356),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(net790),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(net50),
    .X(net1631));
 sky130_fd_sc_hd__clkbuf_2 hold1422 (.A(net3858),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(_00641_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(net792),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(net3186),
    .X(net1635));
 sky130_fd_sc_hd__buf_4 hold1426 (.A(net587),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(_00593_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(net588),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(net3244),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net3062),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 hold1430 (.A(net466),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(_00545_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(net467),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(net3248),
    .X(net1643));
 sky130_fd_sc_hd__buf_4 hold1434 (.A(net583),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(_00561_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(net584),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(net3252),
    .X(net1647));
 sky130_fd_sc_hd__buf_4 hold1438 (.A(net575),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(_00529_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net2551),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(net576),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(net3254),
    .X(net1651));
 sky130_fd_sc_hd__buf_4 hold1442 (.A(net506),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(_00658_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(net507),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(net3840),
    .X(net1655));
 sky130_fd_sc_hd__buf_1 hold1446 (.A(net739),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(net75),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(net740),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(_00586_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net2553),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(net741),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(net3458),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(net817),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(net72),
    .X(net1663));
 sky130_fd_sc_hd__buf_2 hold1454 (.A(net818),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(_00597_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(net819),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(net3256),
    .X(net1667));
 sky130_fd_sc_hd__clkbuf_4 hold1458 (.A(net446),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(net3258),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net2555),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(net447),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(net3264),
    .X(net1671));
 sky130_fd_sc_hd__clkbuf_4 hold1462 (.A(net450),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(net3266),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(net451),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(net2252),
    .X(net1675));
 sky130_fd_sc_hd__buf_1 hold1466 (.A(net772),
    .X(net1676));
 sky130_fd_sc_hd__clkbuf_2 hold1467 (.A(net2302),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_00626_),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(net774),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net3054),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(net3618),
    .X(net1680));
 sky130_fd_sc_hd__clkbuf_4 hold1471 (.A(net252),
    .X(net1681));
 sky130_fd_sc_hd__buf_12 hold1472 (.A(net169),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(net3013),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(net735),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(net3304),
    .X(net1685));
 sky130_fd_sc_hd__buf_4 hold1476 (.A(net662),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(_00659_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(net663),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(net3276),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net3058),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_4 hold1480 (.A(net459),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(net3278),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(net460),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(net3316),
    .X(net1693));
 sky130_fd_sc_hd__buf_4 hold1484 (.A(net668),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(net3770),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(net669),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(net1475),
    .X(net1697));
 sky130_fd_sc_hd__buf_1 hold1488 (.A(net826),
    .X(net1698));
 sky130_fd_sc_hd__buf_1 hold1489 (.A(net1908),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net1577),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_00627_),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(net828),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(net3544),
    .X(net1702));
 sky130_fd_sc_hd__buf_1 hold1493 (.A(net757),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(net136),
    .X(net1704));
 sky130_fd_sc_hd__buf_1 hold1495 (.A(net758),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(net3551),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(net759),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(net3288),
    .X(net1708));
 sky130_fd_sc_hd__clkbuf_4 hold1499 (.A(net468),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net2766),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 hold150 (.A(net1579),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(net3290),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(net469),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(net3284),
    .X(net1712));
 sky130_fd_sc_hd__clkbuf_4 hold1503 (.A(net477),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(net3286),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(net478),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(net3292),
    .X(net1716));
 sky130_fd_sc_hd__clkbuf_4 hold1507 (.A(net475),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(net3294),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(net476),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net1581),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(net3324),
    .X(net1720));
 sky130_fd_sc_hd__clkbuf_4 hold1511 (.A(net488),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_00618_),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(net489),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(net3318),
    .X(net1724));
 sky130_fd_sc_hd__clkbuf_4 hold1515 (.A(net486),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(net3322),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(net487),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(net3296),
    .X(net1728));
 sky130_fd_sc_hd__clkbuf_4 hold1519 (.A(net484),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net2557),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(net3298),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(net485),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(net3306),
    .X(net1732));
 sky130_fd_sc_hd__clkbuf_4 hold1523 (.A(net498),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(net3308),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(net499),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(net3260),
    .X(net1736));
 sky130_fd_sc_hd__clkbuf_4 hold1527 (.A(net518),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(net3262),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(net519),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net2559),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(net3774),
    .X(net1740));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1531 (.A(net713),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(net124),
    .X(net1742));
 sky130_fd_sc_hd__buf_2 hold1533 (.A(net714),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(net3775),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(net715),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(net3310),
    .X(net1746));
 sky130_fd_sc_hd__buf_4 hold1537 (.A(net492),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(net3314),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(net493),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net2561),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(net2321),
    .X(net1750));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold1541 (.A(net880),
    .X(net1751));
 sky130_fd_sc_hd__clkbuf_2 hold1542 (.A(net2373),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(_00634_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(net882),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(net3208),
    .X(net1755));
 sky130_fd_sc_hd__buf_1 hold1546 (.A(net883),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(net884),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_00554_),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(net885),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net3146),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(net3611),
    .X(net1760));
 sky130_fd_sc_hd__buf_1 hold1551 (.A(net949),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(net71),
    .X(net1762));
 sky130_fd_sc_hd__clkbuf_4 hold1553 (.A(net950),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_00598_),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(net951),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(net3326),
    .X(net1766));
 sky130_fd_sc_hd__clkbuf_4 hold1557 (.A(net496),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(net3328),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(net497),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net1522),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\line_buffer.data_out[17] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(net811),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(net49),
    .X(net1772));
 sky130_fd_sc_hd__buf_1 hold1563 (.A(net3851),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(_00642_),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(net813),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(net3268),
    .X(net1776));
 sky130_fd_sc_hd__buf_4 hold1567 (.A(net532),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(net3270),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(net533),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net3064),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\line_buffer.data_out[26] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(net901),
    .X(net1781));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1572 (.A(net3426),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(_00635_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(net903),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(net3280),
    .X(net1785));
 sky130_fd_sc_hd__clkbuf_4 hold1576 (.A(net512),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(net3282),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(net513),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(net3842),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net1362),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(net865),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(net866),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(_00555_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(net867),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(net3466),
    .X(net1795));
 sky130_fd_sc_hd__buf_2 hold1586 (.A(net386),
    .X(net1796));
 sky130_fd_sc_hd__buf_12 hold1587 (.A(net172),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(net2789),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(net816),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net3074),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(net3272),
    .X(net1800));
 sky130_fd_sc_hd__buf_4 hold1591 (.A(net660),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(net3274),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(net661),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(net3300),
    .X(net1804));
 sky130_fd_sc_hd__clkbuf_4 hold1595 (.A(net479),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(net3302),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(net480),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(net3332),
    .X(net1808));
 sky130_fd_sc_hd__clkbuf_4 hold1599 (.A(net504),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net2743),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net1366),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(net3334),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(net505),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(net3462),
    .X(net1812));
 sky130_fd_sc_hd__buf_4 hold1603 (.A(net681),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_00619_),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(net682),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(net3336),
    .X(net1816));
 sky130_fd_sc_hd__buf_4 hold1607 (.A(net500),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(net3338),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(net501),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net2569),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(net3366),
    .X(net1820));
 sky130_fd_sc_hd__clkbuf_4 hold1611 (.A(net510),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(net3370),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(net511),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(net3372),
    .X(net1824));
 sky130_fd_sc_hd__buf_4 hold1615 (.A(net516),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(_00652_),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(net517),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(net3362),
    .X(net1828));
 sky130_fd_sc_hd__buf_4 hold1619 (.A(net524),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net2571),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_00546_),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(net525),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(net3382),
    .X(net1832));
 sky130_fd_sc_hd__buf_4 hold1623 (.A(net526),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(net3384),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(net527),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(net3358),
    .X(net1836));
 sky130_fd_sc_hd__buf_4 hold1627 (.A(net552),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(net3360),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(net553),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net2573),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(net3354),
    .X(net1840));
 sky130_fd_sc_hd__buf_4 hold1631 (.A(net522),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(net3356),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(net523),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(net3344),
    .X(net1844));
 sky130_fd_sc_hd__buf_4 hold1635 (.A(net542),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(net3348),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(net543),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(net3340),
    .X(net1848));
 sky130_fd_sc_hd__clkbuf_4 hold1639 (.A(net544),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net3068),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(net3342),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(net545),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(net3374),
    .X(net1852));
 sky130_fd_sc_hd__buf_4 hold1643 (.A(net563),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(net3376),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(net564),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(net3402),
    .X(net1856));
 sky130_fd_sc_hd__buf_4 hold1647 (.A(net567),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(net3404),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(net568),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net3072),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(net3386),
    .X(net1860));
 sky130_fd_sc_hd__buf_4 hold1651 (.A(net528),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(_00660_),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(net529),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(net1890),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(net1892),
    .X(net1865));
 sky130_fd_sc_hd__clkbuf_4 hold1656 (.A(_03242_),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(net2871),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(net747),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(net3500),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net2604),
    .X(net376));
 sky130_fd_sc_hd__buf_4 hold1660 (.A(net632),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(net3502),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(net633),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(net3512),
    .X(net1873));
 sky130_fd_sc_hd__clkbuf_4 hold1664 (.A(net239),
    .X(net1874));
 sky130_fd_sc_hd__buf_12 hold1665 (.A(net167),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(net2800),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(net676),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(net3412),
    .X(net1878));
 sky130_fd_sc_hd__buf_4 hold1669 (.A(net581),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net2692),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_00644_),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(net582),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(net3406),
    .X(net1882));
 sky130_fd_sc_hd__buf_4 hold1673 (.A(net579),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(net3700),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(net580),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(net3378),
    .X(net1886));
 sky130_fd_sc_hd__buf_4 hold1677 (.A(net548),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(net3380),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(net549),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net2864),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\control_fsm.weight_write_addr[0] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(net1864),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(net454),
    .X(net1892));
 sky130_fd_sc_hd__clkbuf_4 hold1683 (.A(net1865),
    .X(net1893));
 sky130_fd_sc_hd__buf_1 hold1684 (.A(_03271_),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(_00394_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(net456),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(net3388),
    .X(net1897));
 sky130_fd_sc_hd__buf_4 hold1688 (.A(net546),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(net3392),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net1538),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(net547),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\line_buffer.data_out[9] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(net913),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(net44),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(_00650_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(net915),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(net2996),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(net827),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(net1699),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net1052),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net3082),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(net3547),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(net918),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(net3400),
    .X(net1912));
 sky130_fd_sc_hd__buf_4 hold1703 (.A(net571),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_00433_),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(net572),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(net3414),
    .X(net1916));
 sky130_fd_sc_hd__buf_4 hold1707 (.A(net573),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(net3416),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(net574),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net1374),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(net3398),
    .X(net1920));
 sky130_fd_sc_hd__buf_2 hold1711 (.A(net331),
    .X(net1921));
 sky130_fd_sc_hd__clkbuf_16 hold1712 (.A(net173),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(net2810),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(net822),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(net3097),
    .X(net1925));
 sky130_fd_sc_hd__buf_4 hold1716 (.A(net561),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(net3761),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(net562),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(net3394),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(net3077),
    .X(net382));
 sky130_fd_sc_hd__buf_4 hold1720 (.A(net565),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(net3396),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(net566),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(net3548),
    .X(net1933));
 sky130_fd_sc_hd__buf_4 hold1724 (.A(net670),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(_00602_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(net671),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(net3350),
    .X(net1937));
 sky130_fd_sc_hd__buf_4 hold1728 (.A(net559),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(net3352),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net3080),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(net560),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(net3454),
    .X(net1941));
 sky130_fd_sc_hd__buf_4 hold1732 (.A(net554),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(net3456),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(net555),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(net3464),
    .X(net1945));
 sky130_fd_sc_hd__buf_4 hold1736 (.A(net585),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(_00594_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(net586),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(net3486),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net2609),
    .X(net384));
 sky130_fd_sc_hd__buf_4 hold1740 (.A(net569),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(net3679),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(net570),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(net3408),
    .X(net1953));
 sky130_fd_sc_hd__buf_4 hold1744 (.A(net609),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(net3410),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(net610),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(net3608),
    .X(net1957));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1748 (.A(net988),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(net73),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net2850),
    .X(net385));
 sky130_fd_sc_hd__buf_4 hold1750 (.A(net989),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(_00595_),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(net990),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\line_buffer.data_out[18] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(net862),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(net48),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(net863),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(_00643_),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(net864),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\mac_array.mac[7].mac_unit.b[2] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(net3467),
    .X(net386));
 sky130_fd_sc_hd__buf_4 hold1760 (.A(net611),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(net3428),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(net612),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(net3490),
    .X(net1973));
 sky130_fd_sc_hd__buf_4 hold1764 (.A(net599),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(_00588_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(net600),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(net3787),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\line_buffer.data_out[114] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(net2182),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net2684),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(net3577),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(net969),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(net3431),
    .X(net1982));
 sky130_fd_sc_hd__buf_4 hold1773 (.A(net618),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(net3435),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(net619),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(net3439),
    .X(net1986));
 sky130_fd_sc_hd__buf_4 hold1777 (.A(net694),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(net3443),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(net695),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(net1518),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(net3418),
    .X(net1990));
 sky130_fd_sc_hd__buf_4 hold1781 (.A(net603),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(net3422),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(net604),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(net3498),
    .X(net1994));
 sky130_fd_sc_hd__buf_4 hold1785 (.A(net595),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_00621_),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(net596),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(net3468),
    .X(net1998));
 sky130_fd_sc_hd__buf_4 hold1789 (.A(net620),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_03275_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(net3470),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(net621),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(net3482),
    .X(net2002));
 sky130_fd_sc_hd__buf_4 hold1793 (.A(net589),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(net3484),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(net590),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(net2523),
    .X(net2006));
 sky130_fd_sc_hd__buf_1 hold1797 (.A(net895),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(_06370_),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(_06371_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net2746),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net3389),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(_06377_),
    .X(net2010));
 sky130_fd_sc_hd__clkbuf_2 hold1801 (.A(_06384_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(_06424_),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(net2939),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(net300),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(net3789),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(net956),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net2563),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(net3587),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(net966),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(net3474),
    .X(net2022));
 sky130_fd_sc_hd__buf_4 hold1813 (.A(net593),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(net3476),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(net594),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(net3433),
    .X(net2026));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1817 (.A(net461),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(net3492),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(net3493),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net2565),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(net463),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(net3472),
    .X(net2031));
 sky130_fd_sc_hd__buf_2 hold1822 (.A(net350),
    .X(net2032));
 sky130_fd_sc_hd__buf_12 hold1823 (.A(net170),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(net2877),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(net993),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(net3504),
    .X(net2036));
 sky130_fd_sc_hd__buf_4 hold1827 (.A(net601),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(net3508),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(net602),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net2567),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(net3445),
    .X(net2040));
 sky130_fd_sc_hd__buf_4 hold1831 (.A(net616),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(_00425_),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(net617),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(net3510),
    .X(net2044));
 sky130_fd_sc_hd__buf_4 hold1835 (.A(net591),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(net3690),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(net592),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(net3180),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\line_buffer.data_out[115] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(net3085),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(net2398),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(net3497),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(net1011),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\line_buffer.data_out[97] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(net805),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(net93),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(net806),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(_00562_),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(net807),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\line_buffer.data_out[81] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net1378),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(net886),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(net80),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(net887),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(_00578_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(net888),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(net3583),
    .X(net2065));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1856 (.A(net997),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(net3590),
    .X(net2067));
 sky130_fd_sc_hd__buf_1 hold1858 (.A(net998),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(net3598),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net3537),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(net999),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(net3818),
    .X(net2071));
 sky130_fd_sc_hd__buf_1 hold1862 (.A(net874),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(net115),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(net875),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(_00508_),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(net876),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(net3437),
    .X(net2077));
 sky130_fd_sc_hd__buf_4 hold1868 (.A(net607),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(net3641),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(net2676),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(net608),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(net3526),
    .X(net2081));
 sky130_fd_sc_hd__buf_4 hold1872 (.A(net626),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(net3721),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(net627),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(net3536),
    .X(net2085));
 sky130_fd_sc_hd__buf_2 hold1876 (.A(net396),
    .X(net2086));
 sky130_fd_sc_hd__buf_12 hold1877 (.A(net171),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(net2866),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(net894),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net3200),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(net3524),
    .X(net2090));
 sky130_fd_sc_hd__buf_4 hold1881 (.A(net624),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(_00413_),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(net625),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(net3814),
    .X(net2094));
 sky130_fd_sc_hd__buf_1 hold1885 (.A(net958),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(net186),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(net959),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(_00334_),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(net960),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net1555),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(net3534),
    .X(net2100));
 sky130_fd_sc_hd__buf_4 hold1891 (.A(net630),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(_00653_),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(net631),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(net3809),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(net784),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(net785),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(net3810),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(net786),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(net3538),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net2758),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(net1619),
    .X(net400));
 sky130_fd_sc_hd__buf_4 hold1900 (.A(net642),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(_00580_),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(net643),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(net3516),
    .X(net2113));
 sky130_fd_sc_hd__buf_4 hold1904 (.A(net672),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(net3518),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(net673),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(net3185),
    .X(net2117));
 sky130_fd_sc_hd__clkbuf_2 hold1908 (.A(net973),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(net974),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_03274_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(net3192),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(net975),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(net3478),
    .X(net2122));
 sky130_fd_sc_hd__buf_4 hold1913 (.A(net648),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(net3480),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(net649),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(net2998),
    .X(net2126));
 sky130_fd_sc_hd__clkbuf_2 hold1917 (.A(net850),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(net851),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(net3011),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net1623),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(net852),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(net3514),
    .X(net2131));
 sky130_fd_sc_hd__buf_4 hold1922 (.A(net652),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(net3773),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(net653),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(net3815),
    .X(net2135));
 sky130_fd_sc_hd__buf_1 hold1926 (.A(net910),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(net87),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(net911),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(_00570_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net3092),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(net912),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\mac_array.mac[13].mac_unit.b[0] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(net904),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(net162),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(net905),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(_00417_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(net906),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(net3528),
    .X(net2147));
 sky130_fd_sc_hd__buf_4 hold1938 (.A(net634),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(net3532),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net1390),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(net635),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(net3540),
    .X(net2151));
 sky130_fd_sc_hd__buf_4 hold1942 (.A(net646),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(net3669),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(net647),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\mac_array.mac[10].mac_unit.b[0] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(net889),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(net147),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(net890),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(_00441_),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net3090),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(net891),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\mac_array.mac[15].mac_unit.b[6] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(net727),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(net182),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(net728),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(_00340_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(net729),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(net3605),
    .X(net2167));
 sky130_fd_sc_hd__buf_1 hold1958 (.A(net928),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net1382),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(net929),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(_00571_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(net930),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(net3193),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(net3559),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(net1008),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(net3566),
    .X(net2178));
 sky130_fd_sc_hd__buf_4 hold1969 (.A(net656),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net2593),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(_00549_),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(net657),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(net1978),
    .X(net2182));
 sky130_fd_sc_hd__buf_1 hold1973 (.A(net955),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(net941),
    .X(net2184));
 sky130_fd_sc_hd__buf_1 hold1975 (.A(net2019),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(_00547_),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(net957),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(net3520),
    .X(net2188));
 sky130_fd_sc_hd__buf_4 hold1979 (.A(net636),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net2595),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(net3522),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(net637),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(net3824),
    .X(net2192));
 sky130_fd_sc_hd__buf_1 hold1983 (.A(net946),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(net185),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(net947),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(net3825),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(net948),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(net3550),
    .X(net2198));
 sky130_fd_sc_hd__buf_4 hold1989 (.A(net640),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(net2597),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(net3743),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(net641),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(net3821),
    .X(net2202));
 sky130_fd_sc_hd__buf_1 hold1993 (.A(net802),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(net92),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(net803),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(_00563_),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(net804),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(net3578),
    .X(net2208));
 sky130_fd_sc_hd__buf_4 hold1999 (.A(net654),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net1028),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net1058),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net3203),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(_00550_),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(net655),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(\line_buffer.data_out[82] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(net961),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(net79),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(net962),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(_00579_),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(net963),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(net3861),
    .X(net2218));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2009 (.A(net778),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net1565),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(net144),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(net779),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(_00447_),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(net780),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(net3560),
    .X(net2224));
 sky130_fd_sc_hd__buf_4 hold2015 (.A(net664),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(_00629_),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(net665),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(\mac_array.mac[10].mac_unit.b[3] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(net823),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net1384),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(net146),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(net824),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_00444_),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(net825),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(net3588),
    .X(net2234));
 sky130_fd_sc_hd__buf_4 hold2025 (.A(net666),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(_00614_),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(net667),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(net3564),
    .X(net2238));
 sky130_fd_sc_hd__buf_4 hold2029 (.A(net679),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net3088),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(net3652),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(net680),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(net3592),
    .X(net2242));
 sky130_fd_sc_hd__buf_4 hold2033 (.A(net658),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_00620_),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(net659),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(net3570),
    .X(net2246));
 sky130_fd_sc_hd__buf_4 hold2037 (.A(net699),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(_00557_),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(net700),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net3095),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(net3822),
    .X(net2250));
 sky130_fd_sc_hd__clkbuf_2 hold2041 (.A(net952),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(\line_buffer.data_out[33] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(net3630),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(net954),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(net3871),
    .X(net2255));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2046 (.A(net976),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(net95),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(net977),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2049 (.A(_00556_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net1394),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2050 (.A(net978),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2051 (.A(net3596),
    .X(net2261));
 sky130_fd_sc_hd__buf_4 hold2052 (.A(net690),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2053 (.A(_00645_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2054 (.A(net691),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2055 (.A(\line_buffer.data_out[92] ),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2056 (.A(net832),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2057 (.A(net84),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2058 (.A(net833),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2059 (.A(_00573_),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net2645),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2060 (.A(net834),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2061 (.A(net3603),
    .X(net2271));
 sky130_fd_sc_hd__buf_4 hold2062 (.A(net692),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2063 (.A(_00581_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2064 (.A(net693),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2065 (.A(net3552),
    .X(net2275));
 sky130_fd_sc_hd__buf_1 hold2066 (.A(net685),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2067 (.A(net3561),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2068 (.A(net3562),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2069 (.A(net687),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net2648),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2070 (.A(net3022),
    .X(net2280));
 sky130_fd_sc_hd__buf_1 hold2071 (.A(net716),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2072 (.A(net3036),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2073 (.A(net3042),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2074 (.A(net718),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2075 (.A(net2599),
    .X(net2285));
 sky130_fd_sc_hd__clkbuf_4 hold2076 (.A(net2601),
    .X(net2286));
 sky130_fd_sc_hd__buf_12 hold2077 (.A(net176),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2078 (.A(net2831),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2079 (.A(net777),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net2405),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2080 (.A(net3872),
    .X(net2290));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2081 (.A(net799),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2082 (.A(net85),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2083 (.A(net800),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2084 (.A(_00572_),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2085 (.A(net801),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2086 (.A(\mac_array.mac[6].mac_unit.b[2] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2087 (.A(net3235),
    .X(net2297));
 sky130_fd_sc_hd__buf_1 hold2088 (.A(net3236),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2089 (.A(net3237),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net1600),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2090 (.A(net789),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2091 (.A(net3182),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2092 (.A(net773),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2093 (.A(net1677),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2094 (.A(net3614),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2095 (.A(net783),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2096 (.A(net3594),
    .X(net2306));
 sky130_fd_sc_hd__buf_4 hold2097 (.A(net683),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2098 (.A(net3750),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2099 (.A(net684),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net2761),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net2949),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2100 (.A(net3606),
    .X(net2310));
 sky130_fd_sc_hd__buf_4 hold2101 (.A(net688),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2102 (.A(_00596_),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2103 (.A(net689),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2104 (.A(net3830),
    .X(net2314));
 sky130_fd_sc_hd__buf_1 hold2105 (.A(net706),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2106 (.A(net110),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2107 (.A(net707),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2108 (.A(net3831),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2109 (.A(net708),
    .X(net2319));
 sky130_fd_sc_hd__buf_4 hold211 (.A(net2951),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2110 (.A(net3224),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2111 (.A(\line_buffer.data_out[25] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2113 (.A(net3620),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2114 (.A(net1005),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2115 (.A(net3621),
    .X(net2325));
 sky130_fd_sc_hd__buf_2 hold2116 (.A(net329),
    .X(net2326));
 sky130_fd_sc_hd__buf_12 hold2117 (.A(net168),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2118 (.A(net2840),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2119 (.A(net873),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net2953),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2120 (.A(net3069),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2121 (.A(net808),
    .X(net2331));
 sky130_fd_sc_hd__clkbuf_4 hold2123 (.A(net809),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2124 (.A(net3151),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2125 (.A(net810),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2126 (.A(net2854),
    .X(net2336));
 sky130_fd_sc_hd__clkbuf_2 hold2127 (.A(net925),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2129 (.A(net926),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net3106),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2130 (.A(net2858),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2131 (.A(net927),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2132 (.A(net3626),
    .X(net2342));
 sky130_fd_sc_hd__buf_1 hold2133 (.A(net841),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2134 (.A(net150),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2135 (.A(net842),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2136 (.A(_00437_),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2137 (.A(net843),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2138 (.A(net3828),
    .X(net2348));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2139 (.A(net994),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net3108),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2140 (.A(net149),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2141 (.A(net995),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2142 (.A(net3829),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2143 (.A(net996),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2144 (.A(net3823),
    .X(net2354));
 sky130_fd_sc_hd__buf_1 hold2145 (.A(net922),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2146 (.A(net102),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2147 (.A(net923),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2148 (.A(_00533_),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2149 (.A(net924),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net2702),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2150 (.A(\mac_array.mac[5].mac_unit.b[2] ),
    .X(net2360));
 sky130_fd_sc_hd__clkbuf_2 hold2151 (.A(net934),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2152 (.A(net126),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2153 (.A(net935),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2154 (.A(net3860),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2155 (.A(net936),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2156 (.A(net3616),
    .X(net2366));
 sky130_fd_sc_hd__clkbuf_4 hold2157 (.A(net241),
    .X(net2367));
 sky130_fd_sc_hd__buf_12 hold2158 (.A(net166),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2159 (.A(net2770),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net2705),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2160 (.A(net753),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2161 (.A(net3782),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2163 (.A(net881),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2164 (.A(net3636),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2165 (.A(net798),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2166 (.A(\mac_array.mac[4].mac_unit.b[0] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2167 (.A(net835),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2168 (.A(net123),
    .X(net2378));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2169 (.A(net3868),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net3118),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2170 (.A(net3869),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2171 (.A(net837),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2172 (.A(net3844),
    .X(net2382));
 sky130_fd_sc_hd__buf_1 hold2173 (.A(net931),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2174 (.A(net47),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2175 (.A(net932),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2176 (.A(_00646_),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2177 (.A(net933),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2178 (.A(net3241),
    .X(net2388));
 sky130_fd_sc_hd__clkbuf_2 hold2179 (.A(net721),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net3120),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2180 (.A(net3246),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2181 (.A(net3311),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2182 (.A(net723),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2183 (.A(net3168),
    .X(net2393));
 sky130_fd_sc_hd__clkbuf_2 hold2184 (.A(net943),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2185 (.A(net3174),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2186 (.A(net3175),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2187 (.A(net945),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2188 (.A(net2049),
    .X(net2398));
 sky130_fd_sc_hd__buf_1 hold2189 (.A(net940),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(net3110),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2190 (.A(\mac_array.mac[0].mac_unit.b[0] ),
    .X(net2400));
 sky130_fd_sc_hd__clkbuf_2 hold2191 (.A(net2184),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2192 (.A(_00548_),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2193 (.A(net942),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2194 (.A(\control_fsm.weight_write_addr[1] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2195 (.A(net1598),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2196 (.A(net418),
    .X(net2406));
 sky130_fd_sc_hd__clkbuf_2 hold2197 (.A(net1599),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2198 (.A(_03240_),
    .X(net2408));
 sky130_fd_sc_hd__clkbuf_4 hold2199 (.A(net32),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net2753),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net3112),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2200 (.A(net2529),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2201 (.A(net897),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2202 (.A(\mac_array.mac[12].mac_unit.b[6] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2203 (.A(net769),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2204 (.A(net155),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2205 (.A(net770),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2206 (.A(_00431_),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2207 (.A(net771),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2208 (.A(\line_buffer.data_out[29] ),
    .X(net2418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2209 (.A(net829),
    .X(net2419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net2650),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2210 (.A(net52),
    .X(net2420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2211 (.A(net830),
    .X(net2421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2212 (.A(_00638_),
    .X(net2422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2213 (.A(net831),
    .X(net2423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2214 (.A(net3783),
    .X(net2424));
 sky130_fd_sc_hd__buf_1 hold2215 (.A(net838),
    .X(net2425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2216 (.A(net108),
    .X(net2426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2217 (.A(net839),
    .X(net2427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2218 (.A(_00522_),
    .X(net2428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2219 (.A(net840),
    .X(net2429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net2653),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2220 (.A(\mac_array.mac[0].mac_unit.b[3] ),
    .X(net2430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2221 (.A(net766),
    .X(net2431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2222 (.A(net107),
    .X(net2432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2223 (.A(net767),
    .X(net2433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2224 (.A(_00524_),
    .X(net2434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2225 (.A(net768),
    .X(net2435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2226 (.A(net3319),
    .X(net2436));
 sky130_fd_sc_hd__buf_1 hold2227 (.A(net844),
    .X(net2437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2228 (.A(net845),
    .X(net2438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2229 (.A(_00613_),
    .X(net2439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net3114),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2230 (.A(net846),
    .X(net2440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2231 (.A(net2874),
    .X(net2441));
 sky130_fd_sc_hd__clkbuf_2 hold2232 (.A(net1000),
    .X(net2442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2233 (.A(net2995),
    .X(net2443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2234 (.A(_00612_),
    .X(net2444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2235 (.A(net1002),
    .X(net2445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2236 (.A(net3747),
    .X(net2446));
 sky130_fd_sc_hd__clkbuf_2 hold2237 (.A(net736),
    .X(net2447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2238 (.A(net106),
    .X(net2448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2239 (.A(net737),
    .X(net2449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net3116),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2240 (.A(_00525_),
    .X(net2450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2241 (.A(net738),
    .X(net2451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2242 (.A(net3580),
    .X(net2452));
 sky130_fd_sc_hd__buf_1 hold2243 (.A(net853),
    .X(net2453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2244 (.A(net42),
    .X(net2454));
 sky130_fd_sc_hd__clkbuf_2 hold2245 (.A(net854),
    .X(net2455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2246 (.A(_00654_),
    .X(net2456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2247 (.A(net855),
    .X(net2457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2248 (.A(net3494),
    .X(net2458));
 sky130_fd_sc_hd__clkbuf_2 hold2249 (.A(net742),
    .X(net2459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net2720),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2250 (.A(net3530),
    .X(net2460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2251 (.A(net3542),
    .X(net2461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2252 (.A(net744),
    .X(net2462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2253 (.A(net3210),
    .X(net2463));
 sky130_fd_sc_hd__clkbuf_2 hold2254 (.A(net979),
    .X(net2464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2255 (.A(net3219),
    .X(net2465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2256 (.A(net3220),
    .X(net2466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2257 (.A(net981),
    .X(net2467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2258 (.A(net3834),
    .X(net2468));
 sky130_fd_sc_hd__buf_1 hold2259 (.A(net919),
    .X(net2469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(net2723),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2260 (.A(net78),
    .X(net2470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2261 (.A(net920),
    .X(net2471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2262 (.A(_00582_),
    .X(net2472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2263 (.A(net921),
    .X(net2473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2264 (.A(net3624),
    .X(net2474));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2265 (.A(net793),
    .X(net2475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2266 (.A(net111),
    .X(net2476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2267 (.A(net794),
    .X(net2477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2268 (.A(_00517_),
    .X(net2478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2269 (.A(net795),
    .X(net2479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net3122),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2270 (.A(net3798),
    .X(net2480));
 sky130_fd_sc_hd__buf_1 hold2271 (.A(net868),
    .X(net2481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2272 (.A(net112),
    .X(net2482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2273 (.A(net869),
    .X(net2483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2274 (.A(_00516_),
    .X(net2484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2275 (.A(net870),
    .X(net2485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2276 (.A(net3644),
    .X(net2486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2277 (.A(net754),
    .X(net2487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2278 (.A(net40),
    .X(net2488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2279 (.A(net755),
    .X(net2489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net1430),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2280 (.A(_00661_),
    .X(net2490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2281 (.A(net756),
    .X(net2491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2282 (.A(net3833),
    .X(net2492));
 sky130_fd_sc_hd__buf_1 hold2283 (.A(net898),
    .X(net2493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2284 (.A(net39),
    .X(net2494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2285 (.A(net899),
    .X(net2495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2286 (.A(_00662_),
    .X(net2496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2287 (.A(net900),
    .X(net2497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2288 (.A(net3734),
    .X(net2498));
 sky130_fd_sc_hd__buf_1 hold2289 (.A(net907),
    .X(net2499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net2812),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2290 (.A(net137),
    .X(net2500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2291 (.A(net908),
    .X(net2501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2292 (.A(_00459_),
    .X(net2502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2293 (.A(net909),
    .X(net2503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2294 (.A(\mac_array.mac[12].mac_unit.b[7] ),
    .X(net2504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2295 (.A(net847),
    .X(net2505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2296 (.A(net154),
    .X(net2506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2297 (.A(net848),
    .X(net2507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2298 (.A(_00432_),
    .X(net2508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2299 (.A(net849),
    .X(net2509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net1064),
    .X(net233));
 sky130_fd_sc_hd__buf_4 hold230 (.A(net2814),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2300 (.A(net3820),
    .X(net2510));
 sky130_fd_sc_hd__buf_1 hold2301 (.A(net970),
    .X(net2511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2302 (.A(net57),
    .X(net2512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2303 (.A(net971),
    .X(net2513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2304 (.A(_00630_),
    .X(net2514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2305 (.A(net972),
    .X(net2515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2306 (.A(net2583),
    .X(net2516));
 sky130_fd_sc_hd__buf_1 hold2307 (.A(net985),
    .X(net2517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2308 (.A(net2847),
    .X(net2518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2309 (.A(_00628_),
    .X(net2519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net2816),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2310 (.A(net987),
    .X(net2520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2311 (.A(net2859),
    .X(net2521));
 sky130_fd_sc_hd__buf_1 hold2312 (.A(net859),
    .X(net2522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2313 (.A(net3645),
    .X(net2523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2314 (.A(net860),
    .X(net2524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2315 (.A(net2861),
    .X(net2525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2316 (.A(net861),
    .X(net2526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2317 (.A(net3795),
    .X(net2527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2318 (.A(net982),
    .X(net2528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2319 (.A(_00521_),
    .X(net2529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net1437),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2320 (.A(net983),
    .X(net2530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2321 (.A(net3796),
    .X(net2531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2322 (.A(net984),
    .X(net2532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2323 (.A(\mac_array.mac[8].mac_unit.b[1] ),
    .X(net2533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2324 (.A(net748),
    .X(net2534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2325 (.A(net138),
    .X(net2535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2326 (.A(net749),
    .X(net2536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2327 (.A(_00458_),
    .X(net2537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2328 (.A(net750),
    .X(net2538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2329 (.A(\mac_array.mac[12].mac_unit.b[1] ),
    .X(net2539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(net3128),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2330 (.A(net763),
    .X(net2540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2331 (.A(net158),
    .X(net2541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2332 (.A(net764),
    .X(net2542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2333 (.A(_00426_),
    .X(net2543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2334 (.A(net765),
    .X(net2544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2335 (.A(\result[10][1] ),
    .X(net2545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2336 (.A(net347),
    .X(net2546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2337 (.A(_05774_),
    .X(net2547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2338 (.A(net348),
    .X(net2548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2339 (.A(net3453),
    .X(net2549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net2600),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2340 (.A(net349),
    .X(net2550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2341 (.A(\result[0][3] ),
    .X(net2551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2342 (.A(net354),
    .X(net2552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2343 (.A(_06428_),
    .X(net2553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2344 (.A(net355),
    .X(net2554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2345 (.A(net3104),
    .X(net2555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2346 (.A(net356),
    .X(net2556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2347 (.A(\result[10][0] ),
    .X(net2557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2348 (.A(net362),
    .X(net2558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2349 (.A(_05777_),
    .X(net2559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net2660),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2350 (.A(net363),
    .X(net2560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2351 (.A(net3222),
    .X(net2561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2352 (.A(net364),
    .X(net2562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2353 (.A(\result[10][4] ),
    .X(net2563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2354 (.A(net391),
    .X(net2564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2355 (.A(_05768_),
    .X(net2565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2356 (.A(net392),
    .X(net2566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2357 (.A(_00378_),
    .X(net2567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2358 (.A(net393),
    .X(net2568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2359 (.A(\result[11][1] ),
    .X(net2569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net3257),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2360 (.A(net371),
    .X(net2570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2361 (.A(_03233_),
    .X(net2571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2362 (.A(net372),
    .X(net2572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2363 (.A(_00538_),
    .X(net2573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2364 (.A(net373),
    .X(net2574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2365 (.A(\line_buffer.data_out[100] ),
    .X(net2575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2366 (.A(net937),
    .X(net2576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2367 (.A(net90),
    .X(net2577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2368 (.A(net938),
    .X(net2578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2369 (.A(_00565_),
    .X(net2579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net3259),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2370 (.A(net939),
    .X(net2580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2371 (.A(net3647),
    .X(net2581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2372 (.A(net856),
    .X(net2582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2373 (.A(\line_buffer.data_out[35] ),
    .X(net2583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2374 (.A(net857),
    .X(net2584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2375 (.A(_00566_),
    .X(net2585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2376 (.A(net858),
    .X(net2586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2377 (.A(\line_buffer.data_out[99] ),
    .X(net2587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2378 (.A(net877),
    .X(net2588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2379 (.A(net91),
    .X(net2589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(net2627),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2380 (.A(net878),
    .X(net2590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2381 (.A(_00564_),
    .X(net2591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2382 (.A(net879),
    .X(net2592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2383 (.A(\result[11][4] ),
    .X(net2593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2384 (.A(net407),
    .X(net2594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2385 (.A(_03227_),
    .X(net2595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2386 (.A(net408),
    .X(net2596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2387 (.A(_00541_),
    .X(net2597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2388 (.A(net409),
    .X(net2598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2389 (.A(\control_fsm.line_data[5] ),
    .X(net2599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net2630),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2390 (.A(net2285),
    .X(net2600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2391 (.A(net444),
    .X(net2601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2392 (.A(_00391_),
    .X(net2602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2393 (.A(\control_fsm.line_data[4] ),
    .X(net2603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2394 (.A(net1012),
    .X(net2604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2395 (.A(net376),
    .X(net2605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2396 (.A(net1013),
    .X(net2606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2397 (.A(_00390_),
    .X(net2607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2398 (.A(\control_fsm.line_data[3] ),
    .X(net2608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2399 (.A(net1016),
    .X(net2609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net2756),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(net3265),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2400 (.A(net384),
    .X(net2610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2401 (.A(net1017),
    .X(net2611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2402 (.A(_00389_),
    .X(net2612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2403 (.A(net3656),
    .X(net2613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2404 (.A(net1074),
    .X(net2614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2405 (.A(net235),
    .X(net2615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2406 (.A(net1075),
    .X(net2616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2407 (.A(net3658),
    .X(net2617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2408 (.A(net1076),
    .X(net2618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2409 (.A(net236),
    .X(net2619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net3267),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2410 (.A(net1077),
    .X(net2620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2411 (.A(\result_index[2] ),
    .X(net2621));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold2412 (.A(net301),
    .X(net2622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2413 (.A(_00353_),
    .X(net2623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2414 (.A(net1101),
    .X(net2624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2415 (.A(net302),
    .X(net2625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2416 (.A(net1102),
    .X(net2626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2417 (.A(net25),
    .X(net2627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2418 (.A(net448),
    .X(net2628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2419 (.A(_00345_),
    .X(net2629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net3142),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2420 (.A(net1105),
    .X(net2630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2421 (.A(net449),
    .X(net2631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2422 (.A(net1106),
    .X(net2632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2423 (.A(net2693),
    .X(net2633));
 sky130_fd_sc_hd__buf_4 hold2424 (.A(net704),
    .X(net2634));
 sky130_fd_sc_hd__clkbuf_2 hold2425 (.A(_06437_),
    .X(net2635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2426 (.A(_06439_),
    .X(net2636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2427 (.A(_00354_),
    .X(net2637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2428 (.A(net1185),
    .X(net2638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2429 (.A(net276),
    .X(net2639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net3144),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2430 (.A(net27),
    .X(net2640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2431 (.A(net1097),
    .X(net2641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2432 (.A(_00347_),
    .X(net2642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2433 (.A(net1098),
    .X(net2643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2434 (.A(net297),
    .X(net2644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2435 (.A(net29),
    .X(net2645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2436 (.A(net416),
    .X(net2646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2437 (.A(_00349_),
    .X(net2647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2438 (.A(net1140),
    .X(net2648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2439 (.A(net417),
    .X(net2649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net1891),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2440 (.A(net28),
    .X(net2650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2441 (.A(net431),
    .X(net2651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2442 (.A(_00348_),
    .X(net2652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2443 (.A(net1153),
    .X(net2653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2444 (.A(net432),
    .X(net2654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2445 (.A(\line_buffer.data_out[125] ),
    .X(net2655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2446 (.A(net1121),
    .X(net2656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2447 (.A(net101),
    .X(net2657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2448 (.A(net1122),
    .X(net2658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2449 (.A(_00534_),
    .X(net2659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_03272_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2450 (.A(net1123),
    .X(net2660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2451 (.A(\mac_array.mac[8].mac_unit.b[7] ),
    .X(net2661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2452 (.A(net1146),
    .X(net2662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2453 (.A(net711),
    .X(net2663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2454 (.A(net1147),
    .X(net2664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2455 (.A(_00464_),
    .X(net2665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2456 (.A(net1148),
    .X(net2666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2457 (.A(\line_buffer.data_out[45] ),
    .X(net2667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2458 (.A(net1155),
    .X(net2668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2459 (.A(net709),
    .X(net2669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net1895),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2460 (.A(net1156),
    .X(net2670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2461 (.A(_00622_),
    .X(net2671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2462 (.A(net1157),
    .X(net2672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2463 (.A(net3049),
    .X(net2673));
 sky130_fd_sc_hd__buf_2 hold2464 (.A(net1082),
    .X(net2674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2465 (.A(_00419_),
    .X(net2675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2466 (.A(net1083),
    .X(net2676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2467 (.A(net3047),
    .X(net2677));
 sky130_fd_sc_hd__clkbuf_4 hold2468 (.A(net1085),
    .X(net2678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2469 (.A(_00422_),
    .X(net2679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net3132),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2470 (.A(net1086),
    .X(net2680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2471 (.A(net3740),
    .X(net2681));
 sky130_fd_sc_hd__buf_4 hold2472 (.A(net1088),
    .X(net2682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2473 (.A(_00418_),
    .X(net2683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2474 (.A(net1089),
    .X(net2684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2475 (.A(net3695),
    .X(net2685));
 sky130_fd_sc_hd__buf_2 hold2476 (.A(net1091),
    .X(net2686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2477 (.A(_00424_),
    .X(net2687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2478 (.A(net1092),
    .X(net2688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2479 (.A(net3694),
    .X(net2689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net1453),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 hold2480 (.A(net1094),
    .X(net2690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2481 (.A(_00637_),
    .X(net2691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2482 (.A(net1095),
    .X(net2692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2483 (.A(\result_index[0] ),
    .X(net2693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2484 (.A(net2633),
    .X(net2694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2485 (.A(_00351_),
    .X(net2695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2486 (.A(net1111),
    .X(net2696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2487 (.A(\result_index[1] ),
    .X(net2697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2488 (.A(net1113),
    .X(net2698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2489 (.A(_00352_),
    .X(net2699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net3277),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2490 (.A(net1115),
    .X(net2700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2491 (.A(net24),
    .X(net2701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2492 (.A(net1129),
    .X(net2702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2493 (.A(net425),
    .X(net2703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2494 (.A(_00344_),
    .X(net2704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2495 (.A(net1131),
    .X(net2705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2496 (.A(net426),
    .X(net2706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2497 (.A(net22),
    .X(net2707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2498 (.A(net1133),
    .X(net2708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2499 (.A(net464),
    .X(net2709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net2614),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net3279),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2500 (.A(_00342_),
    .X(net2710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2501 (.A(net1135),
    .X(net2711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2502 (.A(net465),
    .X(net2712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2503 (.A(net26),
    .X(net2713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2504 (.A(net1142),
    .X(net2714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2505 (.A(net577),
    .X(net2715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2506 (.A(_00346_),
    .X(net2716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2507 (.A(net1144),
    .X(net2717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2508 (.A(net578),
    .X(net2718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2509 (.A(net23),
    .X(net2719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net2026),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2510 (.A(net1125),
    .X(net2720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2511 (.A(net435),
    .X(net2721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2512 (.A(_00343_),
    .X(net2722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2513 (.A(net1127),
    .X(net2723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2514 (.A(net436),
    .X(net2724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2515 (.A(serial_weight_data[5]),
    .X(net2725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2516 (.A(net1026),
    .X(net2726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2517 (.A(net211),
    .X(net2727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2518 (.A(net1027),
    .X(net2728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2519 (.A(_00403_),
    .X(net2729));
 sky130_fd_sc_hd__buf_4 hold252 (.A(net120),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2520 (.A(net1030),
    .X(net2730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2521 (.A(serial_weight_data[3]),
    .X(net2731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2522 (.A(net1032),
    .X(net2732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2523 (.A(net217),
    .X(net2733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2524 (.A(net1033),
    .X(net2734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2525 (.A(_00401_),
    .X(net2735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2526 (.A(net1036),
    .X(net2736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2527 (.A(serial_weight_data[2]),
    .X(net2737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2528 (.A(net1038),
    .X(net2738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2529 (.A(net214),
    .X(net2739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net2029),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2530 (.A(_00400_),
    .X(net2740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2531 (.A(net1042),
    .X(net2741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2532 (.A(serial_weight_data[4]),
    .X(net2742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2533 (.A(net1050),
    .X(net2743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2534 (.A(net226),
    .X(net2744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2535 (.A(_00402_),
    .X(net2745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2536 (.A(net1054),
    .X(net2746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2537 (.A(serial_weight_data[1]),
    .X(net2747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2538 (.A(net1044),
    .X(net2748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2539 (.A(net220),
    .X(net2749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net2708),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2540 (.A(_00399_),
    .X(net2750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2541 (.A(net1048),
    .X(net2751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2542 (.A(serial_weight_data[7]),
    .X(net2752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2543 (.A(net1062),
    .X(net2753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2544 (.A(net232),
    .X(net2754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2545 (.A(_00405_),
    .X(net2755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2546 (.A(net1066),
    .X(net2756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2547 (.A(serial_weight_data[6]),
    .X(net2757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2548 (.A(net1056),
    .X(net2758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2549 (.A(net229),
    .X(net2759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net2711),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2550 (.A(_00404_),
    .X(net2760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2551 (.A(net1060),
    .X(net2761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2552 (.A(serial_weight_data[0]),
    .X(net2762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2553 (.A(net1068),
    .X(net2763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2554 (.A(net223),
    .X(net2764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2555 (.A(_00398_),
    .X(net2765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2556 (.A(net1072),
    .X(net2766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2557 (.A(\mac_array.mac[11].mac_unit.b[7] ),
    .X(net2767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2558 (.A(net751),
    .X(net2768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2559 (.A(net148),
    .X(net2769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net1639),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2560 (.A(_00440_),
    .X(net2770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2561 (.A(net2369),
    .X(net2771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2562 (.A(net3744),
    .X(net2772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2563 (.A(net814),
    .X(net2773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2567 (.A(_01700_),
    .X(net2777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2569 (.A(_03165_),
    .X(net2779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net1641),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2570 (.A(_03166_),
    .X(net2780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2571 (.A(_03174_),
    .X(net2781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2572 (.A(_03236_),
    .X(net2782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2573 (.A(_00537_),
    .X(net2783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2574 (.A(\control_fsm.weight_write_addr[3] ),
    .X(net2784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2575 (.A(net1340),
    .X(net2785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2576 (.A(net325),
    .X(net2786));
 sky130_fd_sc_hd__clkbuf_4 hold2577 (.A(_03253_),
    .X(net2787));
 sky130_fd_sc_hd__clkbuf_4 hold2578 (.A(_03255_),
    .X(net2788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2579 (.A(_00450_),
    .X(net2789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net3289),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2580 (.A(net1798),
    .X(net2790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2581 (.A(net3729),
    .X(net2791));
 sky130_fd_sc_hd__buf_1 hold2582 (.A(net472),
    .X(net2792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2583 (.A(net41),
    .X(net2793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2584 (.A(_00655_),
    .X(net2794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2585 (.A(net1462),
    .X(net2795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2586 (.A(net474),
    .X(net2796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2587 (.A(\mac_array.mac[2].mac_unit.b[6] ),
    .X(net2797));
 sky130_fd_sc_hd__buf_1 hold2588 (.A(net674),
    .X(net2798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2589 (.A(net113),
    .X(net2799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net3291),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2590 (.A(_00511_),
    .X(net2800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2591 (.A(net1876),
    .X(net2801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2592 (.A(\mac_array.mac[13].mac_unit.b[6] ),
    .X(net2802));
 sky130_fd_sc_hd__buf_1 hold2593 (.A(net1163),
    .X(net2803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2594 (.A(net159),
    .X(net2804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2595 (.A(_00423_),
    .X(net2805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2596 (.A(net1165),
    .X(net2806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2597 (.A(\mac_array.mac[2].mac_unit.b[0] ),
    .X(net2807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2598 (.A(net820),
    .X(net2808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2599 (.A(net116),
    .X(net2809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net2618),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net3134),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2600 (.A(_00505_),
    .X(net2810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2601 (.A(net1923),
    .X(net2811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2602 (.A(\line_buffer.data_out[22] ),
    .X(net2812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2603 (.A(net439),
    .X(net2813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2604 (.A(net46),
    .X(net2814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2605 (.A(_00647_),
    .X(net2815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2606 (.A(net1435),
    .X(net2816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2607 (.A(net441),
    .X(net2817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2608 (.A(\mac_array.mac[9].mac_unit.b[0] ),
    .X(net2818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2609 (.A(net1117),
    .X(net2819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net3136),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2610 (.A(net143),
    .X(net2820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2611 (.A(_00449_),
    .X(net2821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2612 (.A(net1119),
    .X(net2822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2613 (.A(\mac_array.mac[9].mac_unit.b[4] ),
    .X(net2823));
 sky130_fd_sc_hd__buf_1 hold2614 (.A(net1167),
    .X(net2824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2615 (.A(net141),
    .X(net2825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2616 (.A(_00453_),
    .X(net2826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2617 (.A(net1169),
    .X(net2827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2618 (.A(\line_buffer.data_out[93] ),
    .X(net2828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2619 (.A(net775),
    .X(net2829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net2791),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2620 (.A(net83),
    .X(net2830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2621 (.A(_00574_),
    .X(net2831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2622 (.A(net2288),
    .X(net2832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2623 (.A(\control_fsm.state[1] ),
    .X(net2833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2624 (.A(net1020),
    .X(net2834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2625 (.A(net243),
    .X(net2835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2626 (.A(_00356_),
    .X(net2836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2627 (.A(net3882),
    .X(net2837));
 sky130_fd_sc_hd__buf_1 hold2628 (.A(net871),
    .X(net2838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2629 (.A(net125),
    .X(net2839));
 sky130_fd_sc_hd__buf_4 hold263 (.A(net2793),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2630 (.A(_00486_),
    .X(net2840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2631 (.A(net2328),
    .X(net2841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2632 (.A(\control_fsm.weight_write_addr[2] ),
    .X(net2842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2633 (.A(net1544),
    .X(net2843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2634 (.A(net335),
    .X(net2844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2635 (.A(\line_buffer.data_out[27] ),
    .X(net2845));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold2636 (.A(net1171),
    .X(net2846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2637 (.A(net986),
    .X(net2847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2638 (.A(net1172),
    .X(net2848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2639 (.A(_00636_),
    .X(net2849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net2795),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2640 (.A(net1173),
    .X(net2850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2641 (.A(net3819),
    .X(net2851));
 sky130_fd_sc_hd__buf_1 hold2642 (.A(net892),
    .X(net2852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2643 (.A(_03143_),
    .X(net2853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2644 (.A(\mac_array.mac[11].mac_unit.b[3] ),
    .X(net2854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2645 (.A(_03172_),
    .X(net2855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2646 (.A(net2336),
    .X(net2856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2647 (.A(_03234_),
    .X(net2857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2648 (.A(_00436_),
    .X(net2858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2649 (.A(\mac_array.mac[12].mac_unit.b[4] ),
    .X(net2859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net3293),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2650 (.A(net2521),
    .X(net2860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2651 (.A(_00429_),
    .X(net2861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2652 (.A(net2525),
    .X(net2862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2653 (.A(net3878),
    .X(net2863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2654 (.A(net1536),
    .X(net2864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2655 (.A(net378),
    .X(net2865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2656 (.A(_00411_),
    .X(net2866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2657 (.A(net2088),
    .X(net2867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2658 (.A(net3870),
    .X(net2868));
 sky130_fd_sc_hd__buf_1 hold2659 (.A(net745),
    .X(net2869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(net3295),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2660 (.A(net114),
    .X(net2870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2661 (.A(_00509_),
    .X(net2871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2662 (.A(net1867),
    .X(net2872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2663 (.A(net3839),
    .X(net2873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2664 (.A(\line_buffer.data_out[51] ),
    .X(net2874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2666 (.A(net992),
    .X(net2876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2667 (.A(_00468_),
    .X(net2877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2668 (.A(net2034),
    .X(net2878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2669 (.A(\result[13][2] ),
    .X(net2879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net3285),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2670 (.A(net1210),
    .X(net2880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2671 (.A(net261),
    .X(net2881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2672 (.A(_00368_),
    .X(net2882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2673 (.A(net1212),
    .X(net2883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2674 (.A(\result[0][1] ),
    .X(net2884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2675 (.A(net1220),
    .X(net2885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2676 (.A(net257),
    .X(net2886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2677 (.A(_00359_),
    .X(net2887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2678 (.A(net1222),
    .X(net2888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2679 (.A(\result[13][1] ),
    .X(net2889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net3287),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2680 (.A(net1224),
    .X(net2890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2681 (.A(net259),
    .X(net2891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2682 (.A(_00367_),
    .X(net2892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2683 (.A(net1226),
    .X(net2893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2684 (.A(\result[0][6] ),
    .X(net2894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2685 (.A(net1150),
    .X(net2895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2686 (.A(net271),
    .X(net2896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2687 (.A(_00364_),
    .X(net2897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2688 (.A(\mac_array.mac[11].mac_unit.b[1] ),
    .X(net2898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2689 (.A(net1240),
    .X(net2899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net3301),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2690 (.A(net269),
    .X(net2900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2691 (.A(_00434_),
    .X(net2901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2692 (.A(net1242),
    .X(net2902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2693 (.A(\result[10][7] ),
    .X(net2903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2694 (.A(net1228),
    .X(net2904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2695 (.A(net263),
    .X(net2905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2696 (.A(\result[0][2] ),
    .X(net2906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2697 (.A(net1236),
    .X(net2907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2698 (.A(net265),
    .X(net2908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2699 (.A(_00360_),
    .X(net2909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net1215),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net3303),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2700 (.A(net1238),
    .X(net2910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2701 (.A(\result[11][7] ),
    .X(net2911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2702 (.A(net1232),
    .X(net2912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2703 (.A(net267),
    .X(net2913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2704 (.A(\result[13][4] ),
    .X(net2914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2705 (.A(net1250),
    .X(net2915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2706 (.A(net279),
    .X(net2916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2707 (.A(_00370_),
    .X(net2917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2708 (.A(net1252),
    .X(net2918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2709 (.A(\result[0][0] ),
    .X(net2919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net1464),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2710 (.A(net1254),
    .X(net2920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2711 (.A(net277),
    .X(net2921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2712 (.A(_00358_),
    .X(net2922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2713 (.A(net1256),
    .X(net2923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2714 (.A(\result[0][4] ),
    .X(net2924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2715 (.A(net1258),
    .X(net2925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2716 (.A(net273),
    .X(net2926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2717 (.A(_00362_),
    .X(net2927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2718 (.A(\result[13][5] ),
    .X(net2928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2719 (.A(net1268),
    .X(net2929));
 sky130_fd_sc_hd__buf_4 hold272 (.A(net1466),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2720 (.A(net283),
    .X(net2930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2721 (.A(_00371_),
    .X(net2931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2722 (.A(\result[13][6] ),
    .X(net2932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2723 (.A(net1284),
    .X(net2933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2724 (.A(net291),
    .X(net2934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2725 (.A(_00372_),
    .X(net2935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2726 (.A(\result[0][5] ),
    .X(net2936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2727 (.A(net298),
    .X(net2937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2728 (.A(net295),
    .X(net2938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2729 (.A(_00363_),
    .X(net2939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(net1468),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2730 (.A(\line_buffer.data_out[88] ),
    .X(net2940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2731 (.A(net1276),
    .X(net2941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2733 (.A(net1277),
    .X(net2943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2734 (.A(_00569_),
    .X(net2944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2735 (.A(net1278),
    .X(net2945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2736 (.A(\result[13][7] ),
    .X(net2946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2737 (.A(net1288),
    .X(net2947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2738 (.A(net293),
    .X(net2948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2739 (.A(net3835),
    .X(net2949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net3297),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_2 hold2740 (.A(net420),
    .X(net2950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2741 (.A(net56),
    .X(net2951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2742 (.A(_00631_),
    .X(net2952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2743 (.A(net1404),
    .X(net2953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2744 (.A(net422),
    .X(net2954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2745 (.A(\result[10][6] ),
    .X(net2955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2746 (.A(net1272),
    .X(net2956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2747 (.A(net287),
    .X(net2957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2748 (.A(\line_buffer.data_out[10] ),
    .X(net2958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2749 (.A(net1280),
    .X(net2959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net3299),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2751 (.A(net1281),
    .X(net2961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2752 (.A(_00651_),
    .X(net2962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2753 (.A(net1282),
    .X(net2963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2754 (.A(\line_buffer.data_out[109] ),
    .X(net2964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2755 (.A(net1159),
    .X(net2965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2756 (.A(net719),
    .X(net2966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2757 (.A(_00558_),
    .X(net2967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2758 (.A(net1161),
    .X(net2968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2759 (.A(net3811),
    .X(net2969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net1724),
    .X(net486));
 sky130_fd_sc_hd__buf_1 hold2760 (.A(net1175),
    .X(net2970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2762 (.A(net1176),
    .X(net2972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2763 (.A(_00420_),
    .X(net2973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2764 (.A(net1177),
    .X(net2974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2765 (.A(\line_buffer.data_out[122] ),
    .X(net2975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2766 (.A(net1296),
    .X(net2976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2767 (.A(net1297),
    .X(net2977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2768 (.A(_00531_),
    .X(net2978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2769 (.A(net1298),
    .X(net2979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(net3323),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2770 (.A(\result[11][2] ),
    .X(net2980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2771 (.A(net1300),
    .X(net2981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2772 (.A(net309),
    .X(net2982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2773 (.A(_00539_),
    .X(net2983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2774 (.A(\result[11][3] ),
    .X(net2984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2775 (.A(net1316),
    .X(net2985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2776 (.A(net315),
    .X(net2986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2777 (.A(_00540_),
    .X(net2987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2778 (.A(\result[10][3] ),
    .X(net2988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2779 (.A(net1312),
    .X(net2989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(net3325),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2780 (.A(net311),
    .X(net2990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2781 (.A(_00377_),
    .X(net2991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2782 (.A(\result[10][5] ),
    .X(net2992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2783 (.A(net1292),
    .X(net2993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2784 (.A(net313),
    .X(net2994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2785 (.A(net1001),
    .X(net2995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2786 (.A(\line_buffer.data_out[58] ),
    .X(net2996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2787 (.A(net1907),
    .X(net2997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2788 (.A(\mac_array.mac[15].mac_unit.b[4] ),
    .X(net2998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2789 (.A(\line_buffer.data_out[80] ),
    .X(net2999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net1722),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2790 (.A(net1308),
    .X(net3000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2791 (.A(net2126),
    .X(net3001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2792 (.A(net1309),
    .X(net3002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2793 (.A(_00577_),
    .X(net3003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2794 (.A(net1310),
    .X(net3004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2795 (.A(\result[10][2] ),
    .X(net3005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2796 (.A(net1304),
    .X(net3006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2797 (.A(net305),
    .X(net3007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2798 (.A(_00376_),
    .X(net3008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2799 (.A(\mac_array.mac[13].mac_unit.b[4] ),
    .X(net3009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net1205),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net3167),
    .X(net490));
 sky130_fd_sc_hd__buf_1 hold2800 (.A(net733),
    .X(net3010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2801 (.A(_00338_),
    .X(net3011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2802 (.A(net734),
    .X(net3012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2803 (.A(_00421_),
    .X(net3013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2804 (.A(net1683),
    .X(net3014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2805 (.A(\result[11][6] ),
    .X(net3015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2806 (.A(net1320),
    .X(net3016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2807 (.A(net317),
    .X(net3017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2808 (.A(\result[11][5] ),
    .X(net3018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2809 (.A(net1324),
    .X(net3019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net1515),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2810 (.A(net319),
    .X(net3020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2811 (.A(net2129),
    .X(net3021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2812 (.A(\mac_array.mac[6].mac_unit.b[6] ),
    .X(net3022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2815 (.A(net3879),
    .X(net3025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2816 (.A(net1336),
    .X(net3026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2817 (.A(net327),
    .X(net3027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2818 (.A(\line_buffer.data_out[121] ),
    .X(net3028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net1746),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2821 (.A(net1333),
    .X(net3031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2822 (.A(_00530_),
    .X(net3032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2823 (.A(net1334),
    .X(net3033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2824 (.A(\mac_array.mac[9].mac_unit.b[6] ),
    .X(net3034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2825 (.A(net1328),
    .X(net3035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2826 (.A(net717),
    .X(net3036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2827 (.A(net1329),
    .X(net3037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2828 (.A(_00455_),
    .X(net3038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2829 (.A(net1330),
    .X(net3039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net3315),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2830 (.A(\line_buffer.data_out[30] ),
    .X(net3040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2831 (.A(net1344),
    .X(net3041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2832 (.A(_00479_),
    .X(net3042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2833 (.A(net1345),
    .X(net3043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2834 (.A(_00639_),
    .X(net3044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2835 (.A(net1346),
    .X(net3045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2836 (.A(net339),
    .X(net3046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2837 (.A(\mac_array.mac[13].mac_unit.b[5] ),
    .X(net3047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2838 (.A(net2677),
    .X(net3048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2839 (.A(\mac_array.mac[13].mac_unit.b[2] ),
    .X(net3049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net3234),
    .X(net494));
 sky130_fd_sc_hd__buf_1 hold2840 (.A(net1349),
    .X(net3050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2841 (.A(_00471_),
    .X(net3051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2842 (.A(net1350),
    .X(net3052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2843 (.A(\mac_array.mac[14].mac_unit.b[7] ),
    .X(net3053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2844 (.A(net1352),
    .X(net3054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2845 (.A(net2673),
    .X(net3055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2846 (.A(net1353),
    .X(net3056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2847 (.A(_00416_),
    .X(net3057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2848 (.A(net1354),
    .X(net3058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2849 (.A(\line_buffer.data_out[59] ),
    .X(net3059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net1612),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2850 (.A(net1357),
    .X(net3060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2851 (.A(_00604_),
    .X(net3061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2852 (.A(net1358),
    .X(net3062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2853 (.A(\mac_array.mac[8].mac_unit.b[0] ),
    .X(net3063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2854 (.A(net1360),
    .X(net3064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2855 (.A(net367),
    .X(net3065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2856 (.A(_00457_),
    .X(net3066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2857 (.A(\mac_array.mac[10].mac_unit.b[4] ),
    .X(net3067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2858 (.A(net1368),
    .X(net3068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2859 (.A(\mac_array.mac[6].mac_unit.b[0] ),
    .X(net3069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(net3327),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2860 (.A(net1369),
    .X(net3070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2861 (.A(_00445_),
    .X(net3071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2862 (.A(net1370),
    .X(net3072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2863 (.A(\line_buffer.data_out[123] ),
    .X(net3073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2864 (.A(net1364),
    .X(net3074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2865 (.A(net1365),
    .X(net3075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2866 (.A(\result[13][0] ),
    .X(net3076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2867 (.A(net1187),
    .X(net3077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2868 (.A(net382),
    .X(net3078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2869 (.A(_00366_),
    .X(net3079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net3329),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2870 (.A(net1189),
    .X(net3080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2871 (.A(\control_fsm.line_data[0] ),
    .X(net3081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2872 (.A(net1372),
    .X(net3082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2873 (.A(net380),
    .X(net3083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2874 (.A(\control_fsm.line_data[7] ),
    .X(net3084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2875 (.A(net1376),
    .X(net3085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2876 (.A(net394),
    .X(net3086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2877 (.A(_00560_),
    .X(net3087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2878 (.A(net1386),
    .X(net3088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2879 (.A(net3627),
    .X(net3089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net3307),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2880 (.A(net1380),
    .X(net3090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2881 (.A(net3876),
    .X(net3091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2882 (.A(net1388),
    .X(net3092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2883 (.A(net403),
    .X(net3093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2884 (.A(\line_buffer.data_out[23] ),
    .X(net3094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2885 (.A(net1392),
    .X(net3095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2886 (.A(_00648_),
    .X(net3096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2887 (.A(net3760),
    .X(net3097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2888 (.A(net1925),
    .X(net3098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2889 (.A(_06393_),
    .X(net3099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net3309),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2890 (.A(_06394_),
    .X(net3100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2891 (.A(_06395_),
    .X(net3101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2893 (.A(_06398_),
    .X(net3103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2894 (.A(_00361_),
    .X(net3104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2895 (.A(\line_buffer.data_out[55] ),
    .X(net3105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2896 (.A(net1406),
    .X(net3106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2897 (.A(_00616_),
    .X(net3107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2898 (.A(net1408),
    .X(net3108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2899 (.A(\line_buffer.data_out[47] ),
    .X(net3109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net3513),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net3337),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2900 (.A(net1420),
    .X(net3110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2901 (.A(_00624_),
    .X(net3111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2902 (.A(net1422),
    .X(net3112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2903 (.A(\line_buffer.data_out[31] ),
    .X(net3113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2904 (.A(net1424),
    .X(net3114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2905 (.A(_00640_),
    .X(net3115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2906 (.A(net1426),
    .X(net3116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2907 (.A(\line_buffer.data_out[79] ),
    .X(net3117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2908 (.A(net1410),
    .X(net3118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2909 (.A(_00592_),
    .X(net3119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net3339),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2910 (.A(net1412),
    .X(net3120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2911 (.A(net3680),
    .X(net3121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2912 (.A(net1428),
    .X(net3122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2913 (.A(\line_buffer.data_out[63] ),
    .X(net3123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2916 (.A(net1438),
    .X(net3126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2917 (.A(_00608_),
    .X(net3127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2918 (.A(net1439),
    .X(net3128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2919 (.A(net3797),
    .X(net3129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(net1589),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2920 (.A(net1244),
    .X(net3130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2921 (.A(net3748),
    .X(net3131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2922 (.A(net1451),
    .X(net3132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2923 (.A(\line_buffer.data_out[95] ),
    .X(net3133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2924 (.A(net1455),
    .X(net3134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2925 (.A(_00576_),
    .X(net3135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2926 (.A(net1457),
    .X(net3136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2927 (.A(\line_buffer.data_out[46] ),
    .X(net3137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2928 (.A(net1470),
    .X(net3138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2929 (.A(_00623_),
    .X(net3139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net1591),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2930 (.A(net1472),
    .X(net3140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2931 (.A(\line_buffer.data_out[7] ),
    .X(net3141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2932 (.A(net1447),
    .X(net3142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2933 (.A(_00664_),
    .X(net3143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2934 (.A(net1449),
    .X(net3144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2935 (.A(net3873),
    .X(net3145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2936 (.A(net1459),
    .X(net3146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2937 (.A(net365),
    .X(net3147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(net3333),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2940 (.A(net2333),
    .X(net3150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2941 (.A(_00473_),
    .X(net3151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2942 (.A(net557),
    .X(net3152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2943 (.A(_00607_),
    .X(net3153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2944 (.A(net3736),
    .X(net3154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2945 (.A(net1499),
    .X(net3155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2946 (.A(net30),
    .X(net3156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2947 (.A(net1179),
    .X(net3157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2948 (.A(net638),
    .X(net3158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2949 (.A(_00350_),
    .X(net3159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net3335),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2950 (.A(net3705),
    .X(net3160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2951 (.A(net1491),
    .X(net3161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2952 (.A(net3708),
    .X(net3162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2953 (.A(net1503),
    .X(net3163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2954 (.A(net3781),
    .X(net3164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2955 (.A(net1495),
    .X(net3165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2956 (.A(net3771),
    .X(net3166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2957 (.A(net1513),
    .X(net3167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2958 (.A(\mac_array.mac[4].mac_unit.b[3] ),
    .X(net3168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net3255),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2963 (.A(_05129_),
    .X(net3173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2964 (.A(net944),
    .X(net3174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2965 (.A(_00492_),
    .X(net3175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2966 (.A(_06415_),
    .X(net3176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2967 (.A(_06417_),
    .X(net3177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2968 (.A(_06418_),
    .X(net3178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2969 (.A(_06419_),
    .X(net3179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net1653),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2970 (.A(\mac_array.mac[7].mac_unit.b[0] ),
    .X(net3180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2971 (.A(net2048),
    .X(net3181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2972 (.A(\mac_array.mac[6].mac_unit.b[4] ),
    .X(net3182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2973 (.A(net2301),
    .X(net3183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2974 (.A(_00477_),
    .X(net3184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2975 (.A(\mac_array.mac[15].mac_unit.b[3] ),
    .X(net3185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2976 (.A(net3654),
    .X(net3186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2977 (.A(net1635),
    .X(net3187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2978 (.A(_06059_),
    .X(net3188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2979 (.A(net2117),
    .X(net3189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net3138),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2980 (.A(_06067_),
    .X(net3190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2981 (.A(_00369_),
    .X(net3191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2982 (.A(_00337_),
    .X(net3192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2983 (.A(\mac_array.mac[7].mac_unit.b[1] ),
    .X(net3193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2984 (.A(net2173),
    .X(net3194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2985 (.A(net3735),
    .X(net3195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2986 (.A(net1540),
    .X(net3196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2987 (.A(net3762),
    .X(net3197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2988 (.A(net1549),
    .X(net3198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2989 (.A(net3880),
    .X(net3199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net3140),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2990 (.A(net1553),
    .X(net3200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2991 (.A(net398),
    .X(net3201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2992 (.A(net3877),
    .X(net3202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2993 (.A(net1563),
    .X(net3203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2994 (.A(net410),
    .X(net3204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2995 (.A(net1568),
    .X(net3205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2996 (.A(net3712),
    .X(net3206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2997 (.A(net1573),
    .X(net3207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2998 (.A(\line_buffer.data_out[105] ),
    .X(net3208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2999 (.A(net1755),
    .X(net3209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net2730),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net2806),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net1820),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3000 (.A(\mac_array.mac[3].mac_unit.b[3] ),
    .X(net3210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3001 (.A(_04814_),
    .X(net3211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3002 (.A(_04823_),
    .X(net3212));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold3004 (.A(_04858_),
    .X(net3214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3005 (.A(_05641_),
    .X(net3215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3009 (.A(net980),
    .X(net3219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net3371),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3010 (.A(_00500_),
    .X(net3220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3011 (.A(_05778_),
    .X(net3221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3012 (.A(_00374_),
    .X(net3222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3013 (.A(net3670),
    .X(net3223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3014 (.A(\mac_array.mac[6].mac_unit.b[3] ),
    .X(net3224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3015 (.A(net2320),
    .X(net3225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3016 (.A(net1590),
    .X(net3226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3017 (.A(net3758),
    .X(net3227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net3281),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3020 (.A(net1607),
    .X(net3230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3021 (.A(net3780),
    .X(net3231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3022 (.A(net1602),
    .X(net3232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3023 (.A(net3757),
    .X(net3233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3024 (.A(net1610),
    .X(net3234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3025 (.A(net787),
    .X(net3235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3026 (.A(net788),
    .X(net3236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3027 (.A(_00475_),
    .X(net3237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3028 (.A(net1615),
    .X(net3238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3029 (.A(_00601_),
    .X(net3239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net3283),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3030 (.A(net3681),
    .X(net3240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3031 (.A(\mac_array.mac[4].mac_unit.b[4] ),
    .X(net3241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3033 (.A(net1626),
    .X(net3243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3034 (.A(net3653),
    .X(net3244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3036 (.A(net722),
    .X(net3246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3037 (.A(net1640),
    .X(net3247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3038 (.A(net3706),
    .X(net3248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3039 (.A(net1643),
    .X(net3249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(net2698),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3040 (.A(\control_fsm.next_state[0] ),
    .X(net3250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3041 (.A(net1214),
    .X(net3251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3042 (.A(net3674),
    .X(net3252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3043 (.A(net1647),
    .X(net3253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3044 (.A(net3763),
    .X(net3254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3045 (.A(net1651),
    .X(net3255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3046 (.A(\mac_array.mac[5].mac_unit.b[3] ),
    .X(net3256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3047 (.A(net1667),
    .X(net3257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3048 (.A(_00484_),
    .X(net3258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3049 (.A(net1669),
    .X(net3259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net2700),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3050 (.A(\mac_array.mac[9].mac_unit.b[3] ),
    .X(net3260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3051 (.A(net1736),
    .X(net3261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3052 (.A(_00452_),
    .X(net3262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3053 (.A(net1738),
    .X(net3263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3054 (.A(\mac_array.mac[0].mac_unit.b[6] ),
    .X(net3264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3055 (.A(net1671),
    .X(net3265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3056 (.A(_00527_),
    .X(net3266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3057 (.A(net1673),
    .X(net3267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3058 (.A(\mac_array.mac[9].mac_unit.b[7] ),
    .X(net3268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3059 (.A(net1776),
    .X(net3269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net3373),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3060 (.A(_00456_),
    .X(net3270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3061 (.A(net1778),
    .X(net3271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3062 (.A(\mac_array.mac[9].mac_unit.b[5] ),
    .X(net3272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3063 (.A(net1800),
    .X(net3273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3064 (.A(_00454_),
    .X(net3274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3065 (.A(net1802),
    .X(net3275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3066 (.A(\mac_array.mac[2].mac_unit.b[2] ),
    .X(net3276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3067 (.A(net1689),
    .X(net3277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3068 (.A(_00507_),
    .X(net3278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3069 (.A(net1691),
    .X(net3279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net1826),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3070 (.A(\mac_array.mac[9].mac_unit.b[2] ),
    .X(net3280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3071 (.A(net1785),
    .X(net3281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3072 (.A(_00451_),
    .X(net3282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3073 (.A(net1787),
    .X(net3283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3074 (.A(\mac_array.mac[1].mac_unit.b[1] ),
    .X(net3284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3075 (.A(net1712),
    .X(net3285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3076 (.A(_00514_),
    .X(net3286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3077 (.A(net1714),
    .X(net3287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3078 (.A(\mac_array.mac[0].mac_unit.b[7] ),
    .X(net3288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3079 (.A(net1708),
    .X(net3289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(net3261),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3080 (.A(_00528_),
    .X(net3290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3081 (.A(net1710),
    .X(net3291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3082 (.A(\mac_array.mac[1].mac_unit.b[2] ),
    .X(net3292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3083 (.A(net1716),
    .X(net3293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3084 (.A(_00515_),
    .X(net3294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3085 (.A(net1718),
    .X(net3295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3086 (.A(\mac_array.mac[12].mac_unit.b[2] ),
    .X(net3296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3087 (.A(net1728),
    .X(net3297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3088 (.A(_00427_),
    .X(net3298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3089 (.A(net1730),
    .X(net3299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net3263),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3090 (.A(\mac_array.mac[3].mac_unit.b[1] ),
    .X(net3300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3091 (.A(net1804),
    .X(net3301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3092 (.A(_00498_),
    .X(net3302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3093 (.A(net1806),
    .X(net3303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3094 (.A(net3739),
    .X(net3304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3095 (.A(net1685),
    .X(net3305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3096 (.A(\mac_array.mac[10].mac_unit.b[2] ),
    .X(net3306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3097 (.A(net1732),
    .X(net3307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3098 (.A(_00443_),
    .X(net3308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3099 (.A(net1734),
    .X(net3309));
 sky130_fd_sc_hd__buf_1 hold31 (.A(net3639),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net1614),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3100 (.A(\mac_array.mac[4].mac_unit.b[5] ),
    .X(net3310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3101 (.A(_00493_),
    .X(net3311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3102 (.A(net2391),
    .X(net3312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3103 (.A(net1747),
    .X(net3313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3104 (.A(_00494_),
    .X(net3314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3105 (.A(net1748),
    .X(net3315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3106 (.A(\line_buffer.data_out[74] ),
    .X(net3316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3107 (.A(net1693),
    .X(net3317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3108 (.A(\mac_array.mac[14].mac_unit.b[0] ),
    .X(net3318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3109 (.A(\line_buffer.data_out[52] ),
    .X(net3319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net1616),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3111 (.A(net1725),
    .X(net3321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3112 (.A(_00409_),
    .X(net3322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3113 (.A(net1726),
    .X(net3323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3114 (.A(net3704),
    .X(net3324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3115 (.A(net1720),
    .X(net3325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3116 (.A(\mac_array.mac[2].mac_unit.b[1] ),
    .X(net3326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3117 (.A(net1766),
    .X(net3327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3118 (.A(_00506_),
    .X(net3328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3119 (.A(net1768),
    .X(net3329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net3355),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3120 (.A(\next_state[0] ),
    .X(net3330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3121 (.A(net1204),
    .X(net3331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3122 (.A(\mac_array.mac[4].mac_unit.b[1] ),
    .X(net3332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3123 (.A(net1808),
    .X(net3333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3124 (.A(_00490_),
    .X(net3334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3125 (.A(net1810),
    .X(net3335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3126 (.A(\mac_array.mac[8].mac_unit.b[5] ),
    .X(net3336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3127 (.A(net1816),
    .X(net3337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3128 (.A(_00462_),
    .X(net3338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3129 (.A(net1818),
    .X(net3339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net3357),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3130 (.A(\mac_array.mac[8].mac_unit.b[4] ),
    .X(net3340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3131 (.A(net1848),
    .X(net3341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3132 (.A(_00461_),
    .X(net3342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3133 (.A(net1850),
    .X(net3343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3134 (.A(\mac_array.mac[3].mac_unit.b[5] ),
    .X(net3344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3136 (.A(net2437),
    .X(net3346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3137 (.A(net1845),
    .X(net3347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3138 (.A(_00502_),
    .X(net3348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3139 (.A(net1846),
    .X(net3349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(net1828),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3140 (.A(\mac_array.mac[1].mac_unit.b[5] ),
    .X(net3350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3141 (.A(net1937),
    .X(net3351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3142 (.A(_00518_),
    .X(net3352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3143 (.A(net1939),
    .X(net3353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3144 (.A(\mac_array.mac[12].mac_unit.b[5] ),
    .X(net3354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3145 (.A(net1840),
    .X(net3355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3146 (.A(_00430_),
    .X(net3356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3147 (.A(net1842),
    .X(net3357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3148 (.A(\mac_array.mac[5].mac_unit.b[7] ),
    .X(net3358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3149 (.A(net1836),
    .X(net3359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net1830),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3150 (.A(_00488_),
    .X(net3360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3151 (.A(net1838),
    .X(net3361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3152 (.A(net3685),
    .X(net3362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3153 (.A(\control_fsm.line_write_addr[1] ),
    .X(net3363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3154 (.A(net1517),
    .X(net3364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3155 (.A(net1829),
    .X(net3365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3156 (.A(\mac_array.mac[6].mac_unit.b[5] ),
    .X(net3366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3157 (.A(_03273_),
    .X(net3367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3158 (.A(net1521),
    .X(net3368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3159 (.A(net1821),
    .X(net3369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net3383),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3160 (.A(_00478_),
    .X(net3370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3161 (.A(net1822),
    .X(net3371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3162 (.A(net3642),
    .X(net3372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3163 (.A(net1824),
    .X(net3373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3164 (.A(\mac_array.mac[10].mac_unit.b[7] ),
    .X(net3374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3165 (.A(net1852),
    .X(net3375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3166 (.A(_00448_),
    .X(net3376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3167 (.A(net1854),
    .X(net3377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3168 (.A(\mac_array.mac[0].mac_unit.b[5] ),
    .X(net3378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3169 (.A(net1886),
    .X(net3379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net3385),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3170 (.A(_00526_),
    .X(net3380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3171 (.A(net1888),
    .X(net3381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3172 (.A(\mac_array.mac[14].mac_unit.b[3] ),
    .X(net3382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3173 (.A(net1832),
    .X(net3383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3174 (.A(_00412_),
    .X(net3384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3175 (.A(net1834),
    .X(net3385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3176 (.A(net3759),
    .X(net3386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3177 (.A(net1860),
    .X(net3387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3178 (.A(\mac_array.mac[4].mac_unit.b[7] ),
    .X(net3388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3179 (.A(_00383_),
    .X(net3389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net3387),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3181 (.A(net1898),
    .X(net3391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3182 (.A(_00496_),
    .X(net3392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3183 (.A(net1899),
    .X(net3393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3184 (.A(\mac_array.mac[1].mac_unit.b[7] ),
    .X(net3394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3185 (.A(net1929),
    .X(net3395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3186 (.A(_00520_),
    .X(net3396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3187 (.A(net1931),
    .X(net3397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3188 (.A(net3881),
    .X(net3398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3189 (.A(net1920),
    .X(net3399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net1862),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3190 (.A(net3707),
    .X(net3400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3191 (.A(net1912),
    .X(net3401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3192 (.A(\mac_array.mac[2].mac_unit.b[7] ),
    .X(net3402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3193 (.A(net1856),
    .X(net3403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3194 (.A(_00512_),
    .X(net3404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3195 (.A(net1858),
    .X(net3405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3196 (.A(\line_buffer.data_out[77] ),
    .X(net3406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3197 (.A(net1882),
    .X(net3407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3198 (.A(\mac_array.mac[6].mac_unit.b[1] ),
    .X(net3408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3199 (.A(net1953),
    .X(net3409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net2688),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(net1625),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3200 (.A(_00474_),
    .X(net3410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3201 (.A(net1955),
    .X(net3411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3202 (.A(net3722),
    .X(net3412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3203 (.A(net1878),
    .X(net3413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3204 (.A(\mac_array.mac[14].mac_unit.b[6] ),
    .X(net3414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3205 (.A(net1916),
    .X(net3415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3206 (.A(_00415_),
    .X(net3416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3207 (.A(net1918),
    .X(net3417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3208 (.A(\mac_array.mac[3].mac_unit.b[7] ),
    .X(net3418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net1627),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3211 (.A(net1991),
    .X(net3421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3212 (.A(_00504_),
    .X(net3422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3213 (.A(net1992),
    .X(net3423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3216 (.A(net902),
    .X(net3426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3217 (.A(net1970),
    .X(net3427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3218 (.A(_00467_),
    .X(net3428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3219 (.A(net1971),
    .X(net3429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(net3269),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3220 (.A(net1781),
    .X(net3430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3221 (.A(\mac_array.mac[7].mac_unit.b[4] ),
    .X(net3431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3222 (.A(net1782),
    .X(net3432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3223 (.A(\mac_array.mac[4].mac_unit.b[6] ),
    .X(net3433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3224 (.A(net1983),
    .X(net3434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3225 (.A(_00469_),
    .X(net3435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3226 (.A(net1984),
    .X(net3436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3227 (.A(\mac_array.mac[3].mac_unit.b[0] ),
    .X(net3437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3228 (.A(net2077),
    .X(net3438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3229 (.A(\mac_array.mac[7].mac_unit.b[5] ),
    .X(net3439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net3271),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3232 (.A(net1987),
    .X(net3442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3233 (.A(_00470_),
    .X(net3443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3234 (.A(net1988),
    .X(net3444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3235 (.A(net3667),
    .X(net3445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3236 (.A(net2040),
    .X(net3446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3237 (.A(net1902),
    .X(net3447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net3165),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3240 (.A(_05707_),
    .X(net3450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3241 (.A(_05708_),
    .X(net3451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3242 (.A(_05712_),
    .X(net3452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3243 (.A(_00375_),
    .X(net3453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3244 (.A(\mac_array.mac[15].mac_unit.b[5] ),
    .X(net3454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3245 (.A(net1941),
    .X(net3455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3246 (.A(_00339_),
    .X(net3456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3247 (.A(net1943),
    .X(net3457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3248 (.A(\line_buffer.data_out[68] ),
    .X(net3458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3249 (.A(_01873_),
    .X(net3459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(net1497),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3250 (.A(_01874_),
    .X(net3460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3251 (.A(_03125_),
    .X(net3461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3252 (.A(net3778),
    .X(net3462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3253 (.A(net1812),
    .X(net3463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3254 (.A(net3709),
    .X(net3464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3255 (.A(net1945),
    .X(net3465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3256 (.A(net3843),
    .X(net3466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3257 (.A(net1795),
    .X(net3467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3258 (.A(\mac_array.mac[15].mac_unit.b[7] ),
    .X(net3468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3259 (.A(net1998),
    .X(net3469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net1479),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3260 (.A(_00341_),
    .X(net3470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3261 (.A(net2000),
    .X(net3471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3262 (.A(net3816),
    .X(net3472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3263 (.A(net2031),
    .X(net3473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3264 (.A(\mac_array.mac[6].mac_unit.b[7] ),
    .X(net3474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3265 (.A(net2023),
    .X(net3475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3266 (.A(_00480_),
    .X(net3476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3267 (.A(net2024),
    .X(net3477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3268 (.A(\mac_array.mac[14].mac_unit.b[5] ),
    .X(net3478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3269 (.A(net2122),
    .X(net3479));
 sky130_fd_sc_hd__buf_4 hold327 (.A(net1481),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3270 (.A(_00414_),
    .X(net3480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3271 (.A(net2124),
    .X(net3481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3272 (.A(\mac_array.mac[5].mac_unit.b[4] ),
    .X(net3482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3273 (.A(net2002),
    .X(net3483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3274 (.A(_00485_),
    .X(net3484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3275 (.A(net2004),
    .X(net3485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3276 (.A(net3675),
    .X(net3486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3277 (.A(net1949),
    .X(net3487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3278 (.A(net3617),
    .X(net3488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3279 (.A(net1680),
    .X(net3489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net1483),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3280 (.A(\line_buffer.data_out[75] ),
    .X(net3490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3281 (.A(net1973),
    .X(net3491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3282 (.A(net462),
    .X(net3492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3283 (.A(_00495_),
    .X(net3493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3284 (.A(\mac_array.mac[3].mac_unit.b[4] ),
    .X(net3494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3286 (.A(net1010),
    .X(net3496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3287 (.A(_00465_),
    .X(net3497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3288 (.A(net3688),
    .X(net3498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3289 (.A(net1994),
    .X(net3499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(net1485),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3290 (.A(\mac_array.mac[2].mac_unit.b[5] ),
    .X(net3500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3291 (.A(net1869),
    .X(net3501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3292 (.A(_00510_),
    .X(net3502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3293 (.A(net1871),
    .X(net3503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3294 (.A(\mac_array.mac[7].mac_unit.b[7] ),
    .X(net3504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3297 (.A(net2037),
    .X(net3507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3298 (.A(_00472_),
    .X(net3508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3299 (.A(net2038),
    .X(net3509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net2834),
    .X(net243));
 sky130_fd_sc_hd__buf_4 hold330 (.A(net1487),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3300 (.A(net3689),
    .X(net3510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3301 (.A(net2044),
    .X(net3511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3302 (.A(net3838),
    .X(net3512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3303 (.A(net1873),
    .X(net3513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3304 (.A(net3772),
    .X(net3514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3305 (.A(net2131),
    .X(net3515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3306 (.A(\mac_array.mac[10].mac_unit.b[5] ),
    .X(net3516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3307 (.A(net2113),
    .X(net3517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3308 (.A(_00446_),
    .X(net3518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3309 (.A(net2115),
    .X(net3519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net1489),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3310 (.A(\mac_array.mac[0].mac_unit.b[2] ),
    .X(net3520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3311 (.A(net2188),
    .X(net3521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3312 (.A(_00523_),
    .X(net3522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3313 (.A(net2190),
    .X(net3523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3314 (.A(net3625),
    .X(net3524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3315 (.A(net2090),
    .X(net3525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3316 (.A(\line_buffer.data_out[76] ),
    .X(net3526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3317 (.A(net2081),
    .X(net3527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3318 (.A(\mac_array.mac[4].mac_unit.b[2] ),
    .X(net3528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net1844),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3320 (.A(net743),
    .X(net3530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3321 (.A(net2148),
    .X(net3531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3322 (.A(_00491_),
    .X(net3532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3323 (.A(net2149),
    .X(net3533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3324 (.A(net3649),
    .X(net3534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3325 (.A(net2100),
    .X(net3535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3326 (.A(net3859),
    .X(net3536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3327 (.A(net2085),
    .X(net3537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3328 (.A(net3741),
    .X(net3538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3329 (.A(net2109),
    .X(net3539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(net3349),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3330 (.A(net3668),
    .X(net3540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3331 (.A(net2151),
    .X(net3541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3332 (.A(_00501_),
    .X(net3542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3333 (.A(net2461),
    .X(net3543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3334 (.A(\mac_array.mac[8].mac_unit.b[6] ),
    .X(net3544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3335 (.A(net1702),
    .X(net3545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3336 (.A(net917),
    .X(net3546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3337 (.A(_00603_),
    .X(net3547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3338 (.A(net3662),
    .X(net3548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3339 (.A(net1934),
    .X(net3549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net3341),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3340 (.A(net3742),
    .X(net3550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3341 (.A(_00463_),
    .X(net3551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3342 (.A(\mac_array.mac[3].mac_unit.b[6] ),
    .X(net3552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3343 (.A(net2199),
    .X(net3553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3348 (.A(net1007),
    .X(net3558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3349 (.A(_00466_),
    .X(net3559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net3343),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3350 (.A(net3723),
    .X(net3560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3351 (.A(net686),
    .X(net3561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3352 (.A(_00503_),
    .X(net3562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3353 (.A(net2225),
    .X(net3563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3354 (.A(net3650),
    .X(net3564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3355 (.A(net2238),
    .X(net3565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3356 (.A(net3777),
    .X(net3566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3357 (.A(\line_buffer.data_out[78] ),
    .X(net3567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3359 (.A(net2179),
    .X(net3569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net1897),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3360 (.A(net3784),
    .X(net3570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3361 (.A(net2246),
    .X(net3571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3366 (.A(net968),
    .X(net3576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3367 (.A(_00610_),
    .X(net3577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3368 (.A(net3687),
    .X(net3578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3369 (.A(net482),
    .X(net3579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(net3393),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3370 (.A(\line_buffer.data_out[13] ),
    .X(net3580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3371 (.A(net2209),
    .X(net3581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3372 (.A(net2452),
    .X(net3582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3373 (.A(\mac_array.mac[11].mac_unit.b[2] ),
    .X(net3583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3376 (.A(net965),
    .X(net3586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3377 (.A(_00611_),
    .X(net3587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3378 (.A(net3733),
    .X(net3588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net3379),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3380 (.A(net152),
    .X(net3590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3381 (.A(net2235),
    .X(net3591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3382 (.A(net3738),
    .X(net3592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3383 (.A(net2242),
    .X(net3593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3384 (.A(net3749),
    .X(net3594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3385 (.A(net2306),
    .X(net3595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3386 (.A(net3779),
    .X(net3596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3387 (.A(net2261),
    .X(net3597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3388 (.A(_00435_),
    .X(net3598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3389 (.A(\line_buffer.data_out[111] ),
    .X(net3599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net3381),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3390 (.A(net964),
    .X(net3600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3391 (.A(_02117_),
    .X(net3601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3392 (.A(_05721_),
    .X(net3602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3393 (.A(net3776),
    .X(net3603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3394 (.A(net2271),
    .X(net3604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3395 (.A(net3841),
    .X(net3605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3396 (.A(net3648),
    .X(net3606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3397 (.A(net2310),
    .X(net3607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3398 (.A(net3874),
    .X(net3608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3399 (.A(_03193_),
    .X(net3609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_06474_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net3161),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3400 (.A(_03194_),
    .X(net3610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3401 (.A(\line_buffer.data_out[69] ),
    .X(net3611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3402 (.A(net1760),
    .X(net3612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3403 (.A(net782),
    .X(net3613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3404 (.A(net3184),
    .X(net3614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3405 (.A(\control_fsm.weight_data[7] ),
    .X(net3615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3406 (.A(net3638),
    .X(net3616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3407 (.A(\control_fsm.weight_data[4] ),
    .X(net3617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3408 (.A(net3488),
    .X(net3618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3409 (.A(net1004),
    .X(net3619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(net1493),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3410 (.A(_00476_),
    .X(net3620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3411 (.A(\control_fsm.weight_data[5] ),
    .X(net3621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3412 (.A(net2325),
    .X(net3622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3413 (.A(net2331),
    .X(net3623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3414 (.A(\mac_array.mac[1].mac_unit.b[4] ),
    .X(net3624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3415 (.A(\mac_array.mac[14].mac_unit.b[4] ),
    .X(net3625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3416 (.A(\mac_array.mac[11].mac_unit.b[4] ),
    .X(net3626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3417 (.A(\line_buffer.data_out[39] ),
    .X(net3627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3418 (.A(net1381),
    .X(net3628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3419 (.A(net953),
    .X(net3629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net3359),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3420 (.A(_00605_),
    .X(net3630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3424 (.A(net3438),
    .X(net3634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3425 (.A(net797),
    .X(net3635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3426 (.A(_00606_),
    .X(net3636));
 sky130_fd_sc_hd__buf_1 hold3427 (.A(net2419),
    .X(net3637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3428 (.A(net3615),
    .X(net3638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3429 (.A(net2366),
    .X(net3639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net3361),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3430 (.A(net2078),
    .X(net3640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3431 (.A(_00497_),
    .X(net3641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3432 (.A(\line_buffer.data_out[11] ),
    .X(net3642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3433 (.A(net2528),
    .X(net3643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3434 (.A(\line_buffer.data_out[4] ),
    .X(net3644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3435 (.A(net2400),
    .X(net3645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3436 (.A(net2576),
    .X(net3646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3437 (.A(\line_buffer.data_out[101] ),
    .X(net3647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3438 (.A(\line_buffer.data_out[67] ),
    .X(net3648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3439 (.A(\line_buffer.data_out[12] ),
    .X(net3649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net3455),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3440 (.A(\mac_array.mac[5].mac_unit.b[0] ),
    .X(net3650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3441 (.A(net2588),
    .X(net3651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3442 (.A(_00481_),
    .X(net3652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3443 (.A(\line_buffer.data_out[112] ),
    .X(net3653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3444 (.A(\line_buffer.data_out[64] ),
    .X(net3654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3445 (.A(net2383),
    .X(net3655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3446 (.A(\control_fsm.next_state[2] ),
    .X(net3656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3447 (.A(net2613),
    .X(net3657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3448 (.A(\control_fsm.next_state[1] ),
    .X(net3658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3449 (.A(net2617),
    .X(net3659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net3457),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3450 (.A(net3875),
    .X(net3660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3451 (.A(net1396),
    .X(net3661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3452 (.A(\line_buffer.data_out[57] ),
    .X(net3662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3453 (.A(\line_buffer.data_out[56] ),
    .X(net3663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3454 (.A(net556),
    .X(net3664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3455 (.A(_04659_),
    .X(net3665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3456 (.A(_05741_),
    .X(net3666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3457 (.A(\mac_array.mac[12].mac_unit.b[0] ),
    .X(net3667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3458 (.A(\mac_array.mac[11].mac_unit.b[6] ),
    .X(net3668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3459 (.A(_00439_),
    .X(net3669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net1474),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3460 (.A(\line_buffer.data_out[32] ),
    .X(net3670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3461 (.A(net2142),
    .X(net3671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3462 (.A(_06091_),
    .X(net3672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3463 (.A(_06092_),
    .X(net3673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3464 (.A(\line_buffer.data_out[120] ),
    .X(net3674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3465 (.A(\mac_array.mac[10].mac_unit.b[1] ),
    .X(net3675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3466 (.A(net967),
    .X(net3676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3467 (.A(_06225_),
    .X(net3677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3468 (.A(_06226_),
    .X(net3678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3469 (.A(_00442_),
    .X(net3679));
 sky130_fd_sc_hd__buf_4 hold347 (.A(net66),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3470 (.A(\line_buffer.data_out[15] ),
    .X(net3680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3471 (.A(\line_buffer.data_out[48] ),
    .X(net3681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3472 (.A(net2813),
    .X(net3682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3473 (.A(_03840_),
    .X(net3683));
 sky130_fd_sc_hd__buf_1 hold3474 (.A(_03848_),
    .X(net3684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3475 (.A(\line_buffer.data_out[113] ),
    .X(net3685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3476 (.A(_05583_),
    .X(net3686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3477 (.A(\line_buffer.data_out[117] ),
    .X(net3687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3478 (.A(\line_buffer.data_out[44] ),
    .X(net3688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3479 (.A(\mac_array.mac[15].mac_unit.b[1] ),
    .X(net3689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net1477),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3480 (.A(_00335_),
    .X(net3690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3484 (.A(net3832),
    .X(net3694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3485 (.A(net3817),
    .X(net3695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3488 (.A(net1883),
    .X(net3698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3489 (.A(net1558),
    .X(net3699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net3351),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3490 (.A(_00590_),
    .X(net3700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3491 (.A(_01455_),
    .X(net3701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3492 (.A(_03164_),
    .X(net3702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3493 (.A(_03171_),
    .X(net3703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3494 (.A(\line_buffer.data_out[41] ),
    .X(net3704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3495 (.A(\line_buffer.data_out[71] ),
    .X(net3705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3496 (.A(\line_buffer.data_out[96] ),
    .X(net3706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3497 (.A(\mac_array.mac[11].mac_unit.b[0] ),
    .X(net3707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3498 (.A(\line_buffer.data_out[87] ),
    .X(net3708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3499 (.A(\line_buffer.data_out[65] ),
    .X(net3709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net1195),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(net3353),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3500 (.A(net1003),
    .X(net3710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3501 (.A(_05061_),
    .X(net3711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3502 (.A(\line_buffer.data_out[0] ),
    .X(net3712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3506 (.A(_05579_),
    .X(net3716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3509 (.A(net2082),
    .X(net3719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net3098),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3510 (.A(net2413),
    .X(net3720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3511 (.A(_00589_),
    .X(net3721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3512 (.A(\line_buffer.data_out[19] ),
    .X(net3722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3513 (.A(\line_buffer.data_out[36] ),
    .X(net3723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3514 (.A(net2156),
    .X(net3724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3515 (.A(net2540),
    .X(net3725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3516 (.A(_00945_),
    .X(net3726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3517 (.A(_05845_),
    .X(net3727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3518 (.A(_05846_),
    .X(net3728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3519 (.A(\line_buffer.data_out[14] ),
    .X(net3729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(net1927),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3520 (.A(_04080_),
    .X(net3730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3521 (.A(_05754_),
    .X(net3731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3522 (.A(_05755_),
    .X(net3732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3523 (.A(\line_buffer.data_out[53] ),
    .X(net3733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3524 (.A(\mac_array.mac[8].mac_unit.b[2] ),
    .X(net3734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3525 (.A(\line_buffer.data_out[70] ),
    .X(net3735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3526 (.A(\line_buffer.data_out[119] ),
    .X(net3736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3527 (.A(net796),
    .X(net3737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3528 (.A(\line_buffer.data_out[43] ),
    .X(net3738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3529 (.A(\line_buffer.data_out[2] ),
    .X(net3739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(net3375),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3530 (.A(\mac_array.mac[13].mac_unit.b[1] ),
    .X(net3740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3531 (.A(\line_buffer.data_out[83] ),
    .X(net3741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3532 (.A(\mac_array.mac[3].mac_unit.b[2] ),
    .X(net3742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3533 (.A(_00499_),
    .X(net3743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3534 (.A(\mac_array.mac[9].mac_unit.b[1] ),
    .X(net3744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3535 (.A(_05853_),
    .X(net3745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3536 (.A(\line_buffer.data_out[6] ),
    .X(net3746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3537 (.A(\mac_array.mac[0].mac_unit.b[4] ),
    .X(net3747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3538 (.A(\line_buffer.data_out[127] ),
    .X(net3748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3539 (.A(\mac_array.mac[8].mac_unit.b[3] ),
    .X(net3749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(net3377),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3540 (.A(_00460_),
    .X(net3750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3546 (.A(net1974),
    .X(net3756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3547 (.A(\line_buffer.data_out[40] ),
    .X(net3757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3548 (.A(\line_buffer.data_out[24] ),
    .X(net3758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3549 (.A(\line_buffer.data_out[3] ),
    .X(net3759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net3395),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3550 (.A(\mac_array.mac[1].mac_unit.b[0] ),
    .X(net3760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3551 (.A(_00513_),
    .X(net3761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3552 (.A(\line_buffer.data_out[102] ),
    .X(net3762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3553 (.A(\line_buffer.data_out[1] ),
    .X(net3763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3559 (.A(net1694),
    .X(net3769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(net3397),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3560 (.A(_00587_),
    .X(net3770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3561 (.A(\line_buffer.data_out[118] ),
    .X(net3771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3562 (.A(\mac_array.mac[5].mac_unit.b[1] ),
    .X(net3772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3563 (.A(_00482_),
    .X(net3773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3564 (.A(\mac_array.mac[5].mac_unit.b[6] ),
    .X(net3774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3565 (.A(_00487_),
    .X(net3775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3566 (.A(\line_buffer.data_out[84] ),
    .X(net3776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3567 (.A(\line_buffer.data_out[116] ),
    .X(net3777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3568 (.A(\line_buffer.data_out[42] ),
    .X(net3778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3569 (.A(\line_buffer.data_out[20] ),
    .X(net3779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net3403),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3570 (.A(\line_buffer.data_out[104] ),
    .X(net3780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3571 (.A(\line_buffer.data_out[103] ),
    .X(net3781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3572 (.A(\line_buffer.data_out[61] ),
    .X(net3782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3573 (.A(\mac_array.mac[0].mac_unit.b[1] ),
    .X(net3783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3574 (.A(\line_buffer.data_out[108] ),
    .X(net3784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3576 (.A(net1901),
    .X(net3786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3577 (.A(\line_buffer.data_out[49] ),
    .X(net3787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3578 (.A(\line_buffer.data_out[62] ),
    .X(net3788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3579 (.A(\line_buffer.data_out[50] ),
    .X(net3789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(net3405),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3584 (.A(net45),
    .X(net3794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3585 (.A(\mac_array.mac[12].mac_unit.b[3] ),
    .X(net3795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3586 (.A(_00428_),
    .X(net3796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3587 (.A(net21),
    .X(net3797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3588 (.A(\mac_array.mac[1].mac_unit.b[3] ),
    .X(net3798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3589 (.A(_05625_),
    .X(net3799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(net3487),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3599 (.A(\mac_array.mac[14].mac_unit.b[1] ),
    .X(net3809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net1578),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(net1951),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3600 (.A(_00410_),
    .X(net3810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3601 (.A(\mac_array.mac[13].mac_unit.b[3] ),
    .X(net3811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3602 (.A(_02197_),
    .X(net3812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3603 (.A(_03127_),
    .X(net3813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3604 (.A(\mac_array.mac[15].mac_unit.b[0] ),
    .X(net3814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3605 (.A(\line_buffer.data_out[89] ),
    .X(net3815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3606 (.A(\control_fsm.weight_data[3] ),
    .X(net3816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3607 (.A(\mac_array.mac[13].mac_unit.b[7] ),
    .X(net3817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3608 (.A(\mac_array.mac[2].mac_unit.b[3] ),
    .X(net3818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3609 (.A(\mac_array.mac[14].mac_unit.b[2] ),
    .X(net3819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(net3401),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3610 (.A(\line_buffer.data_out[37] ),
    .X(net3820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3611 (.A(\line_buffer.data_out[98] ),
    .X(net3821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3612 (.A(\line_buffer.data_out[60] ),
    .X(net3822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3613 (.A(\line_buffer.data_out[124] ),
    .X(net3823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3614 (.A(\mac_array.mac[15].mac_unit.b[2] ),
    .X(net3824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3615 (.A(_00336_),
    .X(net3825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3616 (.A(\line_buffer.data_out[126] ),
    .X(net3826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3617 (.A(\line_buffer.data_out[94] ),
    .X(net3827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3618 (.A(\mac_array.mac[11].mac_unit.b[5] ),
    .X(net3828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3619 (.A(_00438_),
    .X(net3829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(net1914),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3620 (.A(\mac_array.mac[1].mac_unit.b[6] ),
    .X(net3830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3621 (.A(_00519_),
    .X(net3831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3622 (.A(\line_buffer.data_out[28] ),
    .X(net3832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3623 (.A(\line_buffer.data_out[5] ),
    .X(net3833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3624 (.A(\line_buffer.data_out[85] ),
    .X(net3834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3625 (.A(\line_buffer.data_out[38] ),
    .X(net3835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3627 (.A(_05722_),
    .X(net3837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3628 (.A(\control_fsm.weight_data[6] ),
    .X(net3838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3629 (.A(\mac_array.mac[7].mac_unit.b[3] ),
    .X(net3839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net3415),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3630 (.A(\line_buffer.data_out[73] ),
    .X(net3840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3631 (.A(\line_buffer.data_out[90] ),
    .X(net3841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3632 (.A(\line_buffer.data_out[106] ),
    .X(net3842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3633 (.A(\control_fsm.weight_data[1] ),
    .X(net3843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3634 (.A(\line_buffer.data_out[21] ),
    .X(net3844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(net3417),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3641 (.A(net812),
    .X(net3851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3648 (.A(net791),
    .X(net3858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3649 (.A(\control_fsm.weight_data[2] ),
    .X(net3859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net3253),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3650 (.A(_00483_),
    .X(net3860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3651 (.A(\mac_array.mac[10].mac_unit.b[6] ),
    .X(net3861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3658 (.A(net836),
    .X(net3868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3659 (.A(_00489_),
    .X(net3869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(net1649),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3660 (.A(\mac_array.mac[2].mac_unit.b[4] ),
    .X(net3870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3661 (.A(\line_buffer.data_out[107] ),
    .X(net3871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3662 (.A(\line_buffer.data_out[91] ),
    .X(net3872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3663 (.A(\control_fsm.line_write_addr[2] ),
    .X(net3873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3664 (.A(\line_buffer.data_out[66] ),
    .X(net3874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3665 (.A(\result[11][0] ),
    .X(net3875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3666 (.A(\control_fsm.line_data[6] ),
    .X(net3876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3667 (.A(\control_fsm.line_data[1] ),
    .X(net3877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3668 (.A(\control_fsm.weight_write_enable ),
    .X(net3878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3669 (.A(\control_fsm.line_write_enable ),
    .X(net3879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net2714),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3670 (.A(\control_fsm.line_data[2] ),
    .X(net3880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3671 (.A(\control_fsm.weight_data[0] ),
    .X(net3881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3672 (.A(\mac_array.mac[5].mac_unit.b[5] ),
    .X(net3882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net2717),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(net3407),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net1200),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(net1884),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net3413),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net1880),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(net3249),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(net1645),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(net3465),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(net1947),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(net3187),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net1637),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(net3483),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net1202),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(net3485),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net3511),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net2046),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(net2022),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(net3477),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(net3499),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net1996),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(net3155),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(net1501),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(net3491),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net3130),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(net1975),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(net2036),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(net3509),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(net1990),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(net3423),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(net3232),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(net1604),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(net3634),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(net2079),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(net3409),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net2738),
    .X(net214));
 sky130_fd_sc_hd__buf_2 hold40 (.A(_00692_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(net3411),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(net1969),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(net3429),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(net1507),
    .X(net613));
 sky130_fd_sc_hd__buf_4 hold404 (.A(net1509),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(net1511),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(net3446),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(net2042),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net1982),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net3436),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net1208),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(net3469),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(net3471),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(net3163),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net1505),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net3525),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(net2092),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(net3527),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(net2083),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(net3196),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(net1542),
    .X(net629));
 sky130_fd_sc_hd__buf_1 hold42 (.A(net3489),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(net3535),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net2102),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(net3501),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(net3503),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(net2147),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(net3533),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(net3521),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net3523),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(net3157),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(net1181),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net2827),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(net2198),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(net2200),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(net3539),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(net2111),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net1606),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net1608),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(net3541),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(net2153),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(net3479),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(net3481),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net1594),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(net3198),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net1551),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net3515),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(net2133),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(net2208),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(net2210),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(net2178),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net2180),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(net3593),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net2244),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_06473_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(net3273),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(net3275),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(net3305),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(net1687),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(net2224),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(net2226),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(net2234),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(net2236),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net3317),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(net1695),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net1218),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(net1933),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net1935),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net3517),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(net3519),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(net2797),
    .X(net674));
 sky130_fd_sc_hd__buf_4 hold465 (.A(net2799),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(net2801),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(net3207),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net1575),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net3565),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net2885),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(net2240),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(net3463),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(net1814),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net3595),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(net2308),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(net2275),
    .X(net685));
 sky130_fd_sc_hd__buf_4 hold476 (.A(net117),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(net2278),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(net3607),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(net2312),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net2888),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(net3597),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(net2263),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(net3604),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(net2273),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(net1986),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net3444),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(net1524),
    .X(net696));
 sky130_fd_sc_hd__buf_4 hold487 (.A(net1526),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(net1528),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(net3571),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net2890),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(net2248),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(net1530),
    .X(net701));
 sky130_fd_sc_hd__buf_4 hold492 (.A(net1532),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(net1534),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(net2694),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(net2696),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net2314),
    .X(net706));
 sky130_fd_sc_hd__buf_4 hold497 (.A(net2316),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net2318),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_1 hold499 (.A(net2668),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net1040),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net2893),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(net2672),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_1 hold501 (.A(net2662),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net2666),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net1740),
    .X(net713));
 sky130_fd_sc_hd__buf_4 hold504 (.A(net1742),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(net1744),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net2280),
    .X(net716));
 sky130_fd_sc_hd__buf_4 hold507 (.A(net127),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net2283),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_1 hold509 (.A(net2965),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net2880),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(net2968),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net2388),
    .X(net721));
 sky130_fd_sc_hd__buf_4 hold512 (.A(net121),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net3312),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net1557),
    .X(net724));
 sky130_fd_sc_hd__buf_4 hold515 (.A(net1559),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net1561),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net2161),
    .X(net727));
 sky130_fd_sc_hd__buf_4 hold518 (.A(net2163),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net2165),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net2883),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net1567),
    .X(net730));
 sky130_fd_sc_hd__buf_4 hold521 (.A(net1569),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(net1571),
    .X(net732));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold523 (.A(net3009),
    .X(net733));
 sky130_fd_sc_hd__buf_4 hold524 (.A(net160),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(net3014),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(net2446),
    .X(net736));
 sky130_fd_sc_hd__buf_4 hold527 (.A(net2448),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net2450),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net1655),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net2904),
    .X(net263));
 sky130_fd_sc_hd__buf_4 hold530 (.A(net1657),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net1659),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(net2458),
    .X(net742));
 sky130_fd_sc_hd__buf_4 hold533 (.A(net118),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net3543),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(net2868),
    .X(net745));
 sky130_fd_sc_hd__buf_4 hold536 (.A(net2870),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net2872),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(net2533),
    .X(net748));
 sky130_fd_sc_hd__buf_4 hold539 (.A(net2535),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net1230),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net2537),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(net2767),
    .X(net751));
 sky130_fd_sc_hd__buf_4 hold542 (.A(net2769),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(net2771),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(net2486),
    .X(net754));
 sky130_fd_sc_hd__buf_4 hold545 (.A(net2488),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net2490),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(net3545),
    .X(net757));
 sky130_fd_sc_hd__buf_4 hold548 (.A(net1704),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(net1706),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net2907),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net1583),
    .X(net760));
 sky130_fd_sc_hd__buf_4 hold551 (.A(net1585),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(net1587),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(net2539),
    .X(net763));
 sky130_fd_sc_hd__buf_4 hold554 (.A(net2541),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(net2543),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(net2430),
    .X(net766));
 sky130_fd_sc_hd__buf_4 hold557 (.A(net2432),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(net2434),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net2412),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net2910),
    .X(net266));
 sky130_fd_sc_hd__buf_4 hold560 (.A(net2414),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(net2416),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(net1675),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 hold563 (.A(net60),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(net1678),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(net2828),
    .X(net775));
 sky130_fd_sc_hd__buf_4 hold566 (.A(net2830),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(net2832),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(net2218),
    .X(net778));
 sky130_fd_sc_hd__buf_4 hold569 (.A(net2220),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net2912),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(net2222),
    .X(net780));
 sky130_fd_sc_hd__buf_2 hold571 (.A(net3183),
    .X(net781));
 sky130_fd_sc_hd__buf_4 hold572 (.A(net128),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(net2304),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(net2104),
    .X(net784));
 sky130_fd_sc_hd__buf_4 hold575 (.A(net165),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(net2107),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(net2296),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_4 hold578 (.A(net130),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(net2299),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net1234),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(net1629),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 hold581 (.A(net1631),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(net1633),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net2474),
    .X(net793));
 sky130_fd_sc_hd__buf_4 hold584 (.A(net2476),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(net2478),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(net2371),
    .X(net796));
 sky130_fd_sc_hd__buf_4 hold587 (.A(net67),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(net2374),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(net2290),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net2899),
    .X(net269));
 sky130_fd_sc_hd__buf_4 hold590 (.A(net2292),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(net2294),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(net2202),
    .X(net802));
 sky130_fd_sc_hd__buf_4 hold593 (.A(net2204),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(net2206),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(net2053),
    .X(net805));
 sky130_fd_sc_hd__buf_4 hold596 (.A(net2055),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(net2057),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(net2330),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 hold599 (.A(net131),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net2741),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net2902),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(net2334),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(net1770),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 hold602 (.A(net1772),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(net1774),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(net2772),
    .X(net814));
 sky130_fd_sc_hd__buf_4 hold605 (.A(net142),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(net2790),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(net1661),
    .X(net817));
 sky130_fd_sc_hd__buf_4 hold608 (.A(net1663),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(net1665),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net2895),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(net2807),
    .X(net820));
 sky130_fd_sc_hd__buf_4 hold611 (.A(net2809),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(net2811),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(net2228),
    .X(net823));
 sky130_fd_sc_hd__buf_4 hold614 (.A(net2230),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(net2232),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(net1697),
    .X(net826));
 sky130_fd_sc_hd__buf_4 hold617 (.A(net59),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(net1700),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(net2418),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net1248),
    .X(net272));
 sky130_fd_sc_hd__buf_4 hold620 (.A(net2420),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(net2422),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(net2265),
    .X(net832));
 sky130_fd_sc_hd__buf_4 hold623 (.A(net2267),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(net2269),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(net2376),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_4 hold626 (.A(net2378),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(net2380),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(net2424),
    .X(net838));
 sky130_fd_sc_hd__buf_4 hold629 (.A(net2426),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net2925),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(net2428),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(net2342),
    .X(net841));
 sky130_fd_sc_hd__buf_4 hold632 (.A(net2344),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(net2346),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(net2436),
    .X(net844));
 sky130_fd_sc_hd__buf_4 hold635 (.A(net62),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(net2439),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(net2504),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_4 hold638 (.A(net2506),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(net2508),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net1260),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(net3001),
    .X(net850));
 sky130_fd_sc_hd__buf_4 hold641 (.A(net183),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(net3021),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(net3582),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 hold644 (.A(net2454),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(net2456),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(net2581),
    .X(net856));
 sky130_fd_sc_hd__buf_4 hold647 (.A(net89),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net2585),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(net2860),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net1183),
    .X(net275));
 sky130_fd_sc_hd__buf_4 hold650 (.A(net156),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(net2862),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(net1963),
    .X(net862));
 sky130_fd_sc_hd__buf_4 hold653 (.A(net1965),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(net1967),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(net1789),
    .X(net865));
 sky130_fd_sc_hd__buf_4 hold656 (.A(net96),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(net1793),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(net2480),
    .X(net868));
 sky130_fd_sc_hd__buf_4 hold659 (.A(net2482),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net2638),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(net2484),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net2837),
    .X(net871));
 sky130_fd_sc_hd__buf_4 hold662 (.A(net2839),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(net2841),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net2071),
    .X(net874));
 sky130_fd_sc_hd__buf_4 hold665 (.A(net2073),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(net2075),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net2587),
    .X(net877));
 sky130_fd_sc_hd__buf_4 hold668 (.A(net2589),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(net2591),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net2920),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net1750),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 hold671 (.A(net55),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(net1753),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net3209),
    .X(net883));
 sky130_fd_sc_hd__buf_4 hold674 (.A(net97),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(net1758),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(net2059),
    .X(net886));
 sky130_fd_sc_hd__buf_4 hold677 (.A(net2061),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net2063),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(net2155),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net2923),
    .X(net278));
 sky130_fd_sc_hd__buf_4 hold680 (.A(net2157),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(net2159),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(net2851),
    .X(net892));
 sky130_fd_sc_hd__buf_4 hold683 (.A(net164),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(net2867),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(net2006),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_8 hold686 (.A(net109),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net2410),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(net2492),
    .X(net898));
 sky130_fd_sc_hd__buf_4 hold689 (.A(net2494),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net2915),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(net2496),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(net1780),
    .X(net901));
 sky130_fd_sc_hd__buf_4 hold692 (.A(net54),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(net1783),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(net2141),
    .X(net904));
 sky130_fd_sc_hd__buf_4 hold695 (.A(net2143),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(net2145),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net2498),
    .X(net907));
 sky130_fd_sc_hd__buf_4 hold698 (.A(net2500),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net2502),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net2732),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net2918),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(net2135),
    .X(net910));
 sky130_fd_sc_hd__buf_4 hold701 (.A(net2137),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(net2139),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(net3786),
    .X(net913));
 sky130_fd_sc_hd__buf_4 hold704 (.A(net1903),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(net1905),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_2 hold706 (.A(net2997),
    .X(net916));
 sky130_fd_sc_hd__buf_4 hold707 (.A(net70),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(net1910),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(net2468),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net1263),
    .X(net281));
 sky130_fd_sc_hd__buf_4 hold710 (.A(net2470),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(net2472),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(net2354),
    .X(net922));
 sky130_fd_sc_hd__buf_4 hold713 (.A(net2356),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net2358),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(net2856),
    .X(net925));
 sky130_fd_sc_hd__buf_4 hold716 (.A(net151),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(net2340),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net2167),
    .X(net928));
 sky130_fd_sc_hd__buf_4 hold719 (.A(net86),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(net1266),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(net2171),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(net2382),
    .X(net931));
 sky130_fd_sc_hd__buf_4 hold722 (.A(net2384),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(net2386),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(net2360),
    .X(net934));
 sky130_fd_sc_hd__buf_4 hold725 (.A(net2362),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(net2364),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(net2575),
    .X(net937));
 sky130_fd_sc_hd__buf_4 hold728 (.A(net2577),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(net2579),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net2929),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(net2050),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_4 hold731 (.A(net98),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(net2402),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(net2393),
    .X(net943));
 sky130_fd_sc_hd__buf_4 hold734 (.A(net122),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(net2396),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(net2192),
    .X(net946));
 sky130_fd_sc_hd__buf_4 hold737 (.A(net2194),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(net2196),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(net3612),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net1270),
    .X(net284));
 sky130_fd_sc_hd__buf_4 hold740 (.A(net1762),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(net1764),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(net2250),
    .X(net952));
 sky130_fd_sc_hd__buf_4 hold743 (.A(net68),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(net2253),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(net1979),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_4 hold746 (.A(net99),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(net2186),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(net2094),
    .X(net958));
 sky130_fd_sc_hd__buf_4 hold749 (.A(net2096),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net2959),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(net2098),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(net2212),
    .X(net961));
 sky130_fd_sc_hd__buf_4 hold752 (.A(net2214),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(net2216),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(net2017),
    .X(net964));
 sky130_fd_sc_hd__buf_4 hold755 (.A(net64),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(net2020),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(net1977),
    .X(net967));
 sky130_fd_sc_hd__buf_4 hold758 (.A(net65),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(net1980),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net2963),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(net2510),
    .X(net970));
 sky130_fd_sc_hd__buf_4 hold761 (.A(net2512),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(net2514),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(net3189),
    .X(net973));
 sky130_fd_sc_hd__buf_4 hold764 (.A(net184),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(net2120),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(net2255),
    .X(net976));
 sky130_fd_sc_hd__buf_4 hold767 (.A(net2257),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net2259),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(net2463),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net2956),
    .X(net287));
 sky130_fd_sc_hd__buf_4 hold770 (.A(net119),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net2466),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(net2527),
    .X(net982));
 sky130_fd_sc_hd__buf_4 hold773 (.A(net157),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(net2531),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(net2516),
    .X(net985));
 sky130_fd_sc_hd__buf_4 hold776 (.A(net58),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(net2519),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(net1957),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_2 hold779 (.A(net1959),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net1274),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(net1961),
    .X(net990));
 sky130_fd_sc_hd__buf_1 hold781 (.A(net2873),
    .X(net991));
 sky130_fd_sc_hd__buf_4 hold782 (.A(net133),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(net2878),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(net2348),
    .X(net994));
 sky130_fd_sc_hd__buf_4 hold785 (.A(net2350),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(net2352),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(net2065),
    .X(net997));
 sky130_fd_sc_hd__buf_4 hold788 (.A(net2067),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(net2069),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net2941),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(net2441),
    .X(net1000));
 sky130_fd_sc_hd__buf_4 hold791 (.A(net63),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(net2444),
    .X(net1002));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold793 (.A(net3225),
    .X(net1003));
 sky130_fd_sc_hd__buf_4 hold794 (.A(net129),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(net2323),
    .X(net1005));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold796 (.A(net3194),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 hold797 (.A(net134),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(net2176),
    .X(net1008));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold799 (.A(net3181),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net1034),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net2945),
    .X(net290));
 sky130_fd_sc_hd__buf_4 hold800 (.A(net135),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(net2051),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(net2603),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_2 hold803 (.A(net2605),
    .X(net1013));
 sky130_fd_sc_hd__buf_12 hold804 (.A(net177),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(net2607),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(net2608),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 hold807 (.A(net2610),
    .X(net1017));
 sky130_fd_sc_hd__buf_12 hold808 (.A(net178),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(net2612),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net2933),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(net2833),
    .X(net1020));
 sky130_fd_sc_hd__buf_2 hold811 (.A(net2835),
    .X(net1021));
 sky130_fd_sc_hd__buf_1 hold812 (.A(_00669_),
    .X(net1022));
 sky130_fd_sc_hd__buf_1 hold813 (.A(net1597),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_16 hold814 (.A(_03267_),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(net2602),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(net2725),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(net2727),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(net16),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(net212),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(net1286),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(net2729),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(net213),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(net2731),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(net2733),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(net14),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(net218),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(net2735),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(net219),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(net2737),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(net2739),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net2947),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(net13),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(net215),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(net2740),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(net216),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(net2747),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(net2749),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(net12),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(net221),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(net2750),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(net222),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net1290),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(net2742),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(net2744),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(net15),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(net227),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(net2745),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net228),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(net2757),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(net2759),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(net17),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(net230),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net2937),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(net2760),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(net231),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(net2752),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(net2754),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(net18),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(net233),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(net2755),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(net234),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(net2762),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(net2764),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_06453_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(net11),
    .X(net1070));
 sky130_fd_sc_hd__buf_1 hold861 (.A(net224),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(net2765),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(net225),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(net3657),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(net2615),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(net3659),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(net2619),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(net3251),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(net1216),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net2643),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(net3331),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(net1206),
    .X(net1081));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold872 (.A(net3055),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(net2675),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(net397),
    .X(net1084));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold875 (.A(net3048),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(net2679),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(net330),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(net2681),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(net2683),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net2936),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(net387),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_2 hold881 (.A(net2685),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(net2687),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(net242),
    .X(net1093));
 sky130_fd_sc_hd__buf_2 hold884 (.A(net2689),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(net2691),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(net377),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(net2640),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(net2642),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(net2644),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net2938),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 hold890 (.A(net1108),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(net2623),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(net2625),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(net1107),
    .X(net1103));
 sky130_fd_sc_hd__buf_1 hold894 (.A(net1109),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(net2629),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(net2631),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\state[0] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(net1103),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(net1100),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net2736),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net2015),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 hold900 (.A(net1104),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(net2695),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(net705),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(net2697),
    .X(net1113));
 sky130_fd_sc_hd__buf_4 hold904 (.A(net514),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(net2699),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net515),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(net2818),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 hold908 (.A(net2820),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(net2821),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net2621),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(net332),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(net2655),
    .X(net1121));
 sky130_fd_sc_hd__buf_4 hold912 (.A(net2657),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(net2659),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(net445),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(net2719),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(net2721),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(net2722),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(net2724),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(net2701),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net2624),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(net2703),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(net2704),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(net2706),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(net2707),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(net2709),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(net2710),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(net2712),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(net1262),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(net1264),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(_06447_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net2976),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(net2647),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(net2649),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(net2713),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(net2715),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(net2716),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(net2718),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(net2661),
    .X(net1146));
 sky130_fd_sc_hd__buf_4 hold937 (.A(net2663),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(net2665),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(net712),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net2979),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(net2894),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net2896),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_06450_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(net2652),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(net2654),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(net2667),
    .X(net1155));
 sky130_fd_sc_hd__buf_4 hold946 (.A(net2669),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(net2671),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(net710),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(net2964),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net3006),
    .X(net305));
 sky130_fd_sc_hd__buf_4 hold950 (.A(net2966),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(net2967),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(net720),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(net2802),
    .X(net1163));
 sky130_fd_sc_hd__buf_4 hold954 (.A(net2804),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(net2805),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net240),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(net2823),
    .X(net1167));
 sky130_fd_sc_hd__buf_4 hold958 (.A(net2825),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(net2826),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net1306),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(net253),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(net2845),
    .X(net1171));
 sky130_fd_sc_hd__buf_4 hold962 (.A(net53),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(net2849),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(net385),
    .X(net1174));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold965 (.A(net2969),
    .X(net1175));
 sky130_fd_sc_hd__buf_4 hold966 (.A(net161),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(net2973),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(net351),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(net3156),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net3000),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(net3158),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(net3159),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(net639),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\result_index[3] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(net275),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(net2637),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(net2639),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(net3076),
    .X(net1187));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold978 (.A(net3078),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(net3079),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net3004),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(net383),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(net3364),
    .X(net1191));
 sky130_fd_sc_hd__buf_1 hold982 (.A(net1519),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(_06470_),
    .X(net1193));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold984 (.A(_06471_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(net2836),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(net245),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(net1593),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_2 hold988 (.A(net1595),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(_03263_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net2981),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_06475_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(net247),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_00357_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(net248),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(net3330),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(net1080),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(net238),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(net1081),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_00333_),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(net251),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 input1 (.A(reset),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(serial_line_valid),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(net1069),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(net1045),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(net1039),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(net2734),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(net1051),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net2728),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(net1057),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(net1063),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(serial_weight_valid),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(serial_line_data[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(start),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input3 (.A(serial_line_data[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(serial_line_data[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(serial_line_data[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(serial_line_data[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(serial_line_data[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(serial_line_data[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(serial_line_data[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_16 output21 (.A(net21),
    .X(done));
 sky130_fd_sc_hd__clkbuf_16 output22 (.A(net22),
    .X(serial_result[0]));
 sky130_fd_sc_hd__clkbuf_16 output23 (.A(net23),
    .X(serial_result[1]));
 sky130_fd_sc_hd__clkbuf_16 output24 (.A(net24),
    .X(serial_result[2]));
 sky130_fd_sc_hd__clkbuf_16 output25 (.A(net25),
    .X(serial_result[3]));
 sky130_fd_sc_hd__clkbuf_16 output26 (.A(net26),
    .X(serial_result[4]));
 sky130_fd_sc_hd__clkbuf_16 output27 (.A(net27),
    .X(serial_result[5]));
 sky130_fd_sc_hd__clkbuf_16 output28 (.A(net28),
    .X(serial_result[6]));
 sky130_fd_sc_hd__clkbuf_16 output29 (.A(net29),
    .X(serial_result[7]));
 sky130_fd_sc_hd__clkbuf_16 output30 (.A(net30),
    .X(serial_result_valid));
 sky130_fd_sc_hd__buf_4 wire31 (.A(_03241_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 wire32 (.A(net2408),
    .X(net32));
 sky130_fd_sc_hd__buf_4 wire33 (.A(_00671_),
    .X(net33));
endmodule


magic
tech sky130A
magscale 1 2
timestamp 1717834355
<< obsli1 >>
rect 1104 2159 162840 157777
<< obsm1 >>
rect 1104 2128 162840 157808
<< metal2 >>
rect 13634 159200 13690 160000
rect 40958 159200 41014 160000
rect 68282 159200 68338 160000
rect 95606 159200 95662 160000
rect 122930 159200 122986 160000
rect 150254 159200 150310 160000
rect 7378 0 7434 800
rect 22282 0 22338 800
rect 37186 0 37242 800
rect 52090 0 52146 800
rect 66994 0 67050 800
rect 81898 0 81954 800
rect 96802 0 96858 800
rect 111706 0 111762 800
rect 126610 0 126666 800
rect 141514 0 141570 800
rect 156418 0 156474 800
<< obsm2 >>
rect 1306 159144 13578 159200
rect 13746 159144 40902 159200
rect 41070 159144 68226 159200
rect 68394 159144 95550 159200
rect 95718 159144 122874 159200
rect 123042 159144 150198 159200
rect 150366 159144 162822 159200
rect 1306 856 162822 159144
rect 1306 734 7322 856
rect 7490 734 22226 856
rect 22394 734 37130 856
rect 37298 734 52034 856
rect 52202 734 66938 856
rect 67106 734 81842 856
rect 82010 734 96746 856
rect 96914 734 111650 856
rect 111818 734 126554 856
rect 126722 734 141458 856
rect 141626 734 156362 856
rect 156530 734 162822 856
<< metal3 >>
rect 0 149336 800 149456
rect 163200 146344 164000 146464
rect 0 129480 800 129600
rect 163200 119688 164000 119808
rect 0 109624 800 109744
rect 163200 93032 164000 93152
rect 0 89768 800 89888
rect 0 69912 800 70032
rect 163200 66376 164000 66496
rect 0 50056 800 50176
rect 163200 39720 164000 39840
rect 0 30200 800 30320
rect 163200 13064 164000 13184
rect 0 10344 800 10464
<< obsm3 >>
rect 800 149536 163200 157793
rect 880 149256 163200 149536
rect 800 146544 163200 149256
rect 800 146264 163120 146544
rect 800 129680 163200 146264
rect 880 129400 163200 129680
rect 800 119888 163200 129400
rect 800 119608 163120 119888
rect 800 109824 163200 119608
rect 880 109544 163200 109824
rect 800 93232 163200 109544
rect 800 92952 163120 93232
rect 800 89968 163200 92952
rect 880 89688 163200 89968
rect 800 70112 163200 89688
rect 880 69832 163200 70112
rect 800 66576 163200 69832
rect 800 66296 163120 66576
rect 800 50256 163200 66296
rect 880 49976 163200 50256
rect 800 39920 163200 49976
rect 800 39640 163120 39920
rect 800 30400 163200 39640
rect 880 30120 163200 30400
rect 800 13264 163200 30120
rect 800 12984 163120 13264
rect 800 10544 163200 12984
rect 880 10264 163200 10544
rect 800 2143 163200 10264
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 46059 2347 50208 142765
rect 50688 2347 65568 142765
rect 66048 2347 80928 142765
rect 81408 2347 96288 142765
rect 96768 2347 111648 142765
rect 112128 2347 112733 142765
<< labels >>
rlabel metal2 s 7378 0 7434 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 done
port 2 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 reset
port 3 nsew signal input
rlabel metal2 s 68282 159200 68338 160000 6 serial_line_data[0]
port 4 nsew signal input
rlabel metal2 s 40958 159200 41014 160000 6 serial_line_data[1]
port 5 nsew signal input
rlabel metal2 s 13634 159200 13690 160000 6 serial_line_data[2]
port 6 nsew signal input
rlabel metal3 s 163200 146344 164000 146464 6 serial_line_data[3]
port 7 nsew signal input
rlabel metal3 s 163200 119688 164000 119808 6 serial_line_data[4]
port 8 nsew signal input
rlabel metal3 s 163200 93032 164000 93152 6 serial_line_data[5]
port 9 nsew signal input
rlabel metal3 s 163200 66376 164000 66496 6 serial_line_data[6]
port 10 nsew signal input
rlabel metal3 s 163200 39720 164000 39840 6 serial_line_data[7]
port 11 nsew signal input
rlabel metal2 s 95606 159200 95662 160000 6 serial_line_valid
port 12 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 serial_result[0]
port 13 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 serial_result[1]
port 14 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 serial_result[2]
port 15 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 serial_result[3]
port 16 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 serial_result[4]
port 17 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 serial_result[5]
port 18 nsew signal output
rlabel metal2 s 150254 159200 150310 160000 6 serial_result[6]
port 19 nsew signal output
rlabel metal2 s 122930 159200 122986 160000 6 serial_result[7]
port 20 nsew signal output
rlabel metal3 s 0 129480 800 129600 6 serial_result_valid
port 21 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 serial_weight_data[0]
port 22 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 serial_weight_data[1]
port 23 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 serial_weight_data[2]
port 24 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 serial_weight_data[3]
port 25 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 serial_weight_data[4]
port 26 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 serial_weight_data[5]
port 27 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 serial_weight_data[6]
port 28 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 serial_weight_data[7]
port 29 nsew signal input
rlabel metal3 s 163200 13064 164000 13184 6 serial_weight_valid
port 30 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 start
port 31 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 33 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 164000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29558240
string GDS_FILE /home/designer01/projects/kws_final_final/openlane/kws_final_final/runs/24_06_08_07_52/results/signoff/CNN_Accelerator_Top.magic.gds
string GDS_START 1015452
<< end >>

